module rom(addr,data);
input [13:0] addr;
output reg [7:0] data;
always @(addr) begin
 case(addr)
 0 : data = 8'h81;
 1 : data = 8'hA0;
 2 : data = 8'h01;
 3 : data = 8'h00;
 4 : data = 8'h73;
 5 : data = 8'h2F;
 6 : data = 8'h20;
 7 : data = 8'h34;
 8 : data = 8'hA1;
 9 : data = 8'h4F;
 10 : data = 8'h63;
 11 : data = 8'h06;
 12 : data = 8'hFF;
 13 : data = 8'h03;
 14 : data = 8'hA5;
 15 : data = 8'h4F;
 16 : data = 8'h63;
 17 : data = 8'h03;
 18 : data = 8'hFF;
 19 : data = 8'h03;
 20 : data = 8'hAD;
 21 : data = 8'h4F;
 22 : data = 8'h63;
 23 : data = 8'h00;
 24 : data = 8'hFF;
 25 : data = 8'h03;
 26 : data = 8'h17;
 27 : data = 8'h0F;
 28 : data = 8'h00;
 29 : data = 8'h80;
 30 : data = 8'h13;
 31 : data = 8'h0F;
 32 : data = 8'h6F;
 33 : data = 8'hFE;
 34 : data = 8'h63;
 35 : data = 8'h03;
 36 : data = 8'h0F;
 37 : data = 8'h00;
 38 : data = 8'h02;
 39 : data = 8'h8F;
 40 : data = 8'h73;
 41 : data = 8'h2F;
 42 : data = 8'h20;
 43 : data = 8'h34;
 44 : data = 8'h63;
 45 : data = 8'h53;
 46 : data = 8'h0F;
 47 : data = 8'h00;
 48 : data = 8'h09;
 49 : data = 8'hA0;
 50 : data = 8'h93;
 51 : data = 8'hE1;
 52 : data = 8'h91;
 53 : data = 8'h53;
 54 : data = 8'h17;
 55 : data = 8'h1F;
 56 : data = 8'h00;
 57 : data = 8'h00;
 58 : data = 8'h23;
 59 : data = 8'h25;
 60 : data = 8'h3F;
 61 : data = 8'hFC;
 62 : data = 8'hE5;
 63 : data = 8'hBF;
 64 : data = 8'h73;
 65 : data = 8'h25;
 66 : data = 8'h40;
 67 : data = 8'hF1;
 68 : data = 8'h01;
 69 : data = 8'hE1;
 70 : data = 8'h97;
 71 : data = 8'h02;
 72 : data = 8'h00;
 73 : data = 8'h00;
 74 : data = 8'h93;
 75 : data = 8'h82;
 76 : data = 8'h22;
 77 : data = 8'h01;
 78 : data = 8'h73;
 79 : data = 8'h90;
 80 : data = 8'h52;
 81 : data = 8'h30;
 82 : data = 8'h73;
 83 : data = 8'h50;
 84 : data = 8'h00;
 85 : data = 8'h18;
 86 : data = 8'h01;
 87 : data = 8'h00;
 88 : data = 8'h97;
 89 : data = 8'h02;
 90 : data = 8'h00;
 91 : data = 8'h00;
 92 : data = 8'h93;
 93 : data = 8'h82;
 94 : data = 8'h82;
 95 : data = 8'h01;
 96 : data = 8'h73;
 97 : data = 8'h90;
 98 : data = 8'h52;
 99 : data = 8'h30;
 100 : data = 8'hFD;
 101 : data = 8'h52;
 102 : data = 8'h73;
 103 : data = 8'h90;
 104 : data = 8'h02;
 105 : data = 8'h3B;
 106 : data = 8'hFD;
 107 : data = 8'h42;
 108 : data = 8'h73;
 109 : data = 8'h90;
 110 : data = 8'h02;
 111 : data = 8'h3A;
 112 : data = 8'h97;
 113 : data = 8'h02;
 114 : data = 8'h00;
 115 : data = 8'h00;
 116 : data = 8'h93;
 117 : data = 8'h82;
 118 : data = 8'h82;
 119 : data = 8'h01;
 120 : data = 8'h73;
 121 : data = 8'h90;
 122 : data = 8'h52;
 123 : data = 8'h30;
 124 : data = 8'h73;
 125 : data = 8'h50;
 126 : data = 8'h20;
 127 : data = 8'h30;
 128 : data = 8'h73;
 129 : data = 8'h50;
 130 : data = 8'h30;
 131 : data = 8'h30;
 132 : data = 8'h73;
 133 : data = 8'h50;
 134 : data = 8'h40;
 135 : data = 8'h30;
 136 : data = 8'h81;
 137 : data = 8'h41;
 138 : data = 8'h97;
 139 : data = 8'h02;
 140 : data = 8'h00;
 141 : data = 8'h00;
 142 : data = 8'h93;
 143 : data = 8'h82;
 144 : data = 8'hA2;
 145 : data = 8'hF7;
 146 : data = 8'h73;
 147 : data = 8'h90;
 148 : data = 8'h52;
 149 : data = 8'h30;
 150 : data = 8'h05;
 151 : data = 8'h45;
 152 : data = 8'h7E;
 153 : data = 8'h05;
 154 : data = 8'h63;
 155 : data = 8'h47;
 156 : data = 8'h05;
 157 : data = 8'h00;
 158 : data = 8'h0F;
 159 : data = 8'h00;
 160 : data = 8'hF0;
 161 : data = 8'h0F;
 162 : data = 8'h85;
 163 : data = 8'h41;
 164 : data = 8'h73;
 165 : data = 8'h00;
 166 : data = 8'h00;
 167 : data = 8'h00;
 168 : data = 8'h97;
 169 : data = 8'h02;
 170 : data = 8'h00;
 171 : data = 8'h80;
 172 : data = 8'h93;
 173 : data = 8'h82;
 174 : data = 8'h82;
 175 : data = 8'hF5;
 176 : data = 8'h63;
 177 : data = 8'h8E;
 178 : data = 8'h02;
 179 : data = 8'h00;
 180 : data = 8'h73;
 181 : data = 8'h90;
 182 : data = 8'h52;
 183 : data = 8'h10;
 184 : data = 8'hB7;
 185 : data = 8'hB2;
 186 : data = 8'h00;
 187 : data = 8'h00;
 188 : data = 8'h93;
 189 : data = 8'h82;
 190 : data = 8'h92;
 191 : data = 8'h10;
 192 : data = 8'h73;
 193 : data = 8'h90;
 194 : data = 8'h22;
 195 : data = 8'h30;
 196 : data = 8'h73;
 197 : data = 8'h23;
 198 : data = 8'h20;
 199 : data = 8'h30;
 200 : data = 8'hE3;
 201 : data = 8'h95;
 202 : data = 8'h62;
 203 : data = 8'hF6;
 204 : data = 8'h73;
 205 : data = 8'h50;
 206 : data = 8'h00;
 207 : data = 8'h30;
 208 : data = 8'h37;
 209 : data = 8'h25;
 210 : data = 8'h00;
 211 : data = 8'h00;
 212 : data = 8'h13;
 213 : data = 8'h05;
 214 : data = 8'h05;
 215 : data = 8'h80;
 216 : data = 8'h73;
 217 : data = 8'h20;
 218 : data = 8'h05;
 219 : data = 8'h30;
 220 : data = 8'h97;
 221 : data = 8'h02;
 222 : data = 8'h00;
 223 : data = 8'h00;
 224 : data = 8'h93;
 225 : data = 8'h82;
 226 : data = 8'h42;
 227 : data = 8'h01;
 228 : data = 8'h73;
 229 : data = 8'h90;
 230 : data = 8'h12;
 231 : data = 8'h34;
 232 : data = 8'h73;
 233 : data = 8'h25;
 234 : data = 8'h40;
 235 : data = 8'hF1;
 236 : data = 8'h73;
 237 : data = 8'h00;
 238 : data = 8'h20;
 239 : data = 8'h30;
 240 : data = 8'h17;
 241 : data = 8'h21;
 242 : data = 8'h00;
 243 : data = 8'h00;
 244 : data = 8'h13;
 245 : data = 8'h01;
 246 : data = 8'h01;
 247 : data = 8'hF1;
 248 : data = 8'h01;
 249 : data = 8'h42;
 250 : data = 8'h81;
 251 : data = 8'h41;
 252 : data = 8'h92;
 253 : data = 8'h91;
 254 : data = 8'h0E;
 255 : data = 8'hC0;
 256 : data = 8'h81;
 257 : data = 8'h44;
 258 : data = 8'h05;
 259 : data = 8'h44;
 260 : data = 8'h26;
 261 : data = 8'h94;
 262 : data = 8'h22;
 263 : data = 8'hC2;
 264 : data = 8'h01;
 265 : data = 8'h46;
 266 : data = 8'h93;
 267 : data = 8'h05;
 268 : data = 8'hF0;
 269 : data = 8'hFF;
 270 : data = 8'hB2;
 271 : data = 8'h95;
 272 : data = 8'h2E;
 273 : data = 8'hC4;
 274 : data = 8'h01;
 275 : data = 8'h47;
 276 : data = 8'hB7;
 277 : data = 8'h86;
 278 : data = 8'h00;
 279 : data = 8'h00;
 280 : data = 8'h93;
 281 : data = 8'h86;
 282 : data = 8'hF6;
 283 : data = 8'hFF;
 284 : data = 8'hBA;
 285 : data = 8'h96;
 286 : data = 8'h36;
 287 : data = 8'hC6;
 288 : data = 8'h01;
 289 : data = 8'h48;
 290 : data = 8'hA1;
 291 : data = 8'h67;
 292 : data = 8'hC2;
 293 : data = 8'h97;
 294 : data = 8'h3E;
 295 : data = 8'hC8;
 296 : data = 8'h17;
 297 : data = 8'h21;
 298 : data = 8'h00;
 299 : data = 8'h00;
 300 : data = 8'h13;
 301 : data = 8'h01;
 302 : data = 8'hC1;
 303 : data = 8'hEE;
 304 : data = 8'h05;
 305 : data = 8'h49;
 306 : data = 8'h81;
 307 : data = 8'h48;
 308 : data = 8'hCA;
 309 : data = 8'h98;
 310 : data = 8'h46;
 311 : data = 8'hC0;
 312 : data = 8'h05;
 313 : data = 8'h4A;
 314 : data = 8'h85;
 315 : data = 8'h49;
 316 : data = 8'hD2;
 317 : data = 8'h99;
 318 : data = 8'h4E;
 319 : data = 8'hC2;
 320 : data = 8'h05;
 321 : data = 8'h4B;
 322 : data = 8'h93;
 323 : data = 8'h0A;
 324 : data = 8'hF0;
 325 : data = 8'hFF;
 326 : data = 8'hDA;
 327 : data = 8'h9A;
 328 : data = 8'h56;
 329 : data = 8'hC4;
 330 : data = 8'h05;
 331 : data = 8'h4C;
 332 : data = 8'hB7;
 333 : data = 8'h8B;
 334 : data = 8'h00;
 335 : data = 8'h00;
 336 : data = 8'h93;
 337 : data = 8'h8B;
 338 : data = 8'hFB;
 339 : data = 8'hFF;
 340 : data = 8'hE2;
 341 : data = 8'h9B;
 342 : data = 8'h5E;
 343 : data = 8'hC6;
 344 : data = 8'h05;
 345 : data = 8'h4D;
 346 : data = 8'hA1;
 347 : data = 8'h6C;
 348 : data = 8'hEA;
 349 : data = 8'h9C;
 350 : data = 8'h66;
 351 : data = 8'hC8;
 352 : data = 8'h17;
 353 : data = 8'h21;
 354 : data = 8'h00;
 355 : data = 8'h00;
 356 : data = 8'h13;
 357 : data = 8'h01;
 358 : data = 8'h81;
 359 : data = 8'hEC;
 360 : data = 8'h13;
 361 : data = 8'h0E;
 362 : data = 8'hF0;
 363 : data = 8'hFF;
 364 : data = 8'h81;
 365 : data = 8'h4D;
 366 : data = 8'hF2;
 367 : data = 8'h9D;
 368 : data = 8'h6E;
 369 : data = 8'hC0;
 370 : data = 8'h13;
 371 : data = 8'h0F;
 372 : data = 8'hF0;
 373 : data = 8'hFF;
 374 : data = 8'h85;
 375 : data = 8'h4E;
 376 : data = 8'hFA;
 377 : data = 8'h9E;
 378 : data = 8'h76;
 379 : data = 8'hC2;
 380 : data = 8'h93;
 381 : data = 8'h01;
 382 : data = 8'hF0;
 383 : data = 8'hFF;
 384 : data = 8'h93;
 385 : data = 8'h0A;
 386 : data = 8'hF0;
 387 : data = 8'hFF;
 388 : data = 8'h8E;
 389 : data = 8'h9A;
 390 : data = 8'h56;
 391 : data = 8'hC4;
 392 : data = 8'h13;
 393 : data = 8'h04;
 394 : data = 8'hF0;
 395 : data = 8'hFF;
 396 : data = 8'h37;
 397 : data = 8'h82;
 398 : data = 8'h00;
 399 : data = 8'h00;
 400 : data = 8'h13;
 401 : data = 8'h02;
 402 : data = 8'hF2;
 403 : data = 8'hFF;
 404 : data = 8'h22;
 405 : data = 8'h92;
 406 : data = 8'h12;
 407 : data = 8'hC6;
 408 : data = 8'h93;
 409 : data = 8'h05;
 410 : data = 8'hF0;
 411 : data = 8'hFF;
 412 : data = 8'hA1;
 413 : data = 8'h64;
 414 : data = 8'hAE;
 415 : data = 8'h94;
 416 : data = 8'h26;
 417 : data = 8'hC8;
 418 : data = 8'h17;
 419 : data = 8'h21;
 420 : data = 8'h00;
 421 : data = 8'h00;
 422 : data = 8'h13;
 423 : data = 8'h01;
 424 : data = 8'hA1;
 425 : data = 8'hE9;
 426 : data = 8'hB7;
 427 : data = 8'h86;
 428 : data = 8'h00;
 429 : data = 8'h00;
 430 : data = 8'h93;
 431 : data = 8'h86;
 432 : data = 8'hF6;
 433 : data = 8'hFF;
 434 : data = 8'h01;
 435 : data = 8'h46;
 436 : data = 8'h36;
 437 : data = 8'h96;
 438 : data = 8'h32;
 439 : data = 8'hC0;
 440 : data = 8'hB7;
 441 : data = 8'h87;
 442 : data = 8'h00;
 443 : data = 8'h00;
 444 : data = 8'h93;
 445 : data = 8'h87;
 446 : data = 8'hF7;
 447 : data = 8'hFF;
 448 : data = 8'h05;
 449 : data = 8'h47;
 450 : data = 8'h3E;
 451 : data = 8'h97;
 452 : data = 8'h3A;
 453 : data = 8'hC2;
 454 : data = 8'hB7;
 455 : data = 8'h88;
 456 : data = 8'h00;
 457 : data = 8'h00;
 458 : data = 8'h93;
 459 : data = 8'h88;
 460 : data = 8'hF8;
 461 : data = 8'hFF;
 462 : data = 8'h13;
 463 : data = 8'h08;
 464 : data = 8'hF0;
 465 : data = 8'hFF;
 466 : data = 8'h46;
 467 : data = 8'h98;
 468 : data = 8'h42;
 469 : data = 8'hC4;
 470 : data = 8'hB7;
 471 : data = 8'h89;
 472 : data = 8'h00;
 473 : data = 8'h00;
 474 : data = 8'h93;
 475 : data = 8'h89;
 476 : data = 8'hF9;
 477 : data = 8'hFF;
 478 : data = 8'h37;
 479 : data = 8'h89;
 480 : data = 8'h00;
 481 : data = 8'h00;
 482 : data = 8'h13;
 483 : data = 8'h09;
 484 : data = 8'hF9;
 485 : data = 8'hFF;
 486 : data = 8'h4E;
 487 : data = 8'h99;
 488 : data = 8'h4A;
 489 : data = 8'hC6;
 490 : data = 8'hB7;
 491 : data = 8'h8A;
 492 : data = 8'h00;
 493 : data = 8'h00;
 494 : data = 8'h93;
 495 : data = 8'h8A;
 496 : data = 8'hFA;
 497 : data = 8'hFF;
 498 : data = 8'h21;
 499 : data = 8'h6A;
 500 : data = 8'h56;
 501 : data = 8'h9A;
 502 : data = 8'h52;
 503 : data = 8'hC8;
 504 : data = 8'h17;
 505 : data = 8'h21;
 506 : data = 8'h00;
 507 : data = 8'h00;
 508 : data = 8'h13;
 509 : data = 8'h01;
 510 : data = 8'h81;
 511 : data = 8'hE5;
 512 : data = 8'hA1;
 513 : data = 8'h6B;
 514 : data = 8'h01;
 515 : data = 8'h4B;
 516 : data = 8'h5E;
 517 : data = 8'h9B;
 518 : data = 8'h5A;
 519 : data = 8'hC0;
 520 : data = 8'hA1;
 521 : data = 8'h6C;
 522 : data = 8'h05;
 523 : data = 8'h4C;
 524 : data = 8'h66;
 525 : data = 8'h9C;
 526 : data = 8'h62;
 527 : data = 8'hC2;
 528 : data = 8'hA1;
 529 : data = 8'h6D;
 530 : data = 8'h13;
 531 : data = 8'h0D;
 532 : data = 8'hF0;
 533 : data = 8'hFF;
 534 : data = 8'h6E;
 535 : data = 8'h9D;
 536 : data = 8'h6A;
 537 : data = 8'hC4;
 538 : data = 8'hA1;
 539 : data = 8'h6E;
 540 : data = 8'h37;
 541 : data = 8'h8E;
 542 : data = 8'h00;
 543 : data = 8'h00;
 544 : data = 8'h13;
 545 : data = 8'h0E;
 546 : data = 8'hFE;
 547 : data = 8'hFF;
 548 : data = 8'h76;
 549 : data = 8'h9E;
 550 : data = 8'h72;
 551 : data = 8'hC6;
 552 : data = 8'hA1;
 553 : data = 8'h6A;
 554 : data = 8'h21;
 555 : data = 8'h6F;
 556 : data = 8'h56;
 557 : data = 8'h9F;
 558 : data = 8'h7A;
 559 : data = 8'hC8;
 560 : data = 8'h0F;
 561 : data = 8'h00;
 562 : data = 8'hF0;
 563 : data = 8'h0F;
 564 : data = 8'h85;
 565 : data = 8'h41;
 566 : data = 8'h73;
 567 : data = 8'h00;
 568 : data = 8'h00;
 569 : data = 8'h00;
 570 : data = 8'h00;
 571 : data = 8'h00;
 572 : data = 8'h00;
 573 : data = 8'h00;
 574 : data = 8'h00;
 575 : data = 8'h00;
 576 : data = 8'h00;
 577 : data = 8'h00;
 578 : data = 8'h00;
 579 : data = 8'h00;
 580 : data = 8'h00;
 581 : data = 8'h00;
 582 : data = 8'h00;
 583 : data = 8'h00;
 584 : data = 8'h00;
 585 : data = 8'h00;
 586 : data = 8'h00;
 587 : data = 8'h00;
 588 : data = 8'h00;
 589 : data = 8'h00;
 590 : data = 8'h00;
 591 : data = 8'h00;
 592 : data = 8'h00;
 593 : data = 8'h00;
 594 : data = 8'h00;
 595 : data = 8'h00;
 596 : data = 8'h00;
 597 : data = 8'h00;
 598 : data = 8'h00;
 599 : data = 8'h00;
 600 : data = 8'h00;
 601 : data = 8'h00;
 602 : data = 8'h00;
 603 : data = 8'h00;
 604 : data = 8'h00;
 605 : data = 8'h00;
 606 : data = 8'h00;
 607 : data = 8'h00;
 608 : data = 8'h00;
 609 : data = 8'h00;
 610 : data = 8'h00;
 611 : data = 8'h00;
 612 : data = 8'h00;
 613 : data = 8'h00;
 614 : data = 8'h00;
 615 : data = 8'h00;
 616 : data = 8'h00;
 617 : data = 8'h00;
 618 : data = 8'h00;
 619 : data = 8'h00;
 620 : data = 8'h00;
 621 : data = 8'h00;
 622 : data = 8'h00;
 623 : data = 8'h00;
 624 : data = 8'h00;
 625 : data = 8'h00;
 626 : data = 8'h00;
 627 : data = 8'h00;
 628 : data = 8'h00;
 629 : data = 8'h00;
 630 : data = 8'h00;
 631 : data = 8'h00;
 632 : data = 8'h00;
 633 : data = 8'h00;
 634 : data = 8'h00;
 635 : data = 8'h00;
 636 : data = 8'h00;
 637 : data = 8'h00;
 638 : data = 8'h00;
 639 : data = 8'h00;
 640 : data = 8'h00;
 641 : data = 8'h00;
 642 : data = 8'h00;
 643 : data = 8'h00;
 644 : data = 8'h00;
 645 : data = 8'h00;
 646 : data = 8'h00;
 647 : data = 8'h00;
 648 : data = 8'h00;
 649 : data = 8'h00;
 650 : data = 8'h00;
 651 : data = 8'h00;
 652 : data = 8'h00;
 653 : data = 8'h00;
 654 : data = 8'h00;
 655 : data = 8'h00;
 656 : data = 8'h00;
 657 : data = 8'h00;
 658 : data = 8'h00;
 659 : data = 8'h00;
 660 : data = 8'h00;
 661 : data = 8'h00;
 662 : data = 8'h00;
 663 : data = 8'h00;
 664 : data = 8'h00;
 665 : data = 8'h00;
 666 : data = 8'h00;
 667 : data = 8'h00;
 668 : data = 8'h00;
 669 : data = 8'h00;
 670 : data = 8'h00;
 671 : data = 8'h00;
 672 : data = 8'h00;
 673 : data = 8'h00;
 674 : data = 8'h00;
 675 : data = 8'h00;
 676 : data = 8'h00;
 677 : data = 8'h00;
 678 : data = 8'h00;
 679 : data = 8'h00;
 680 : data = 8'h00;
 681 : data = 8'h00;
 682 : data = 8'h00;
 683 : data = 8'h00;
 684 : data = 8'h00;
 685 : data = 8'h00;
 686 : data = 8'h00;
 687 : data = 8'h00;
 688 : data = 8'h00;
 689 : data = 8'h00;
 690 : data = 8'h00;
 691 : data = 8'h00;
 692 : data = 8'h00;
 693 : data = 8'h00;
 694 : data = 8'h00;
 695 : data = 8'h00;
 696 : data = 8'h00;
 697 : data = 8'h00;
 698 : data = 8'h00;
 699 : data = 8'h00;
 700 : data = 8'h00;
 701 : data = 8'h00;
 702 : data = 8'h00;
 703 : data = 8'h00;
 704 : data = 8'h00;
 705 : data = 8'h00;
 706 : data = 8'h00;
 707 : data = 8'h00;
 708 : data = 8'h00;
 709 : data = 8'h00;
 710 : data = 8'h00;
 711 : data = 8'h00;
 712 : data = 8'h00;
 713 : data = 8'h00;
 714 : data = 8'h00;
 715 : data = 8'h00;
 716 : data = 8'h00;
 717 : data = 8'h00;
 718 : data = 8'h00;
 719 : data = 8'h00;
 720 : data = 8'h00;
 721 : data = 8'h00;
 722 : data = 8'h00;
 723 : data = 8'h00;
 724 : data = 8'h00;
 725 : data = 8'h00;
 726 : data = 8'h00;
 727 : data = 8'h00;
 728 : data = 8'h00;
 729 : data = 8'h00;
 730 : data = 8'h00;
 731 : data = 8'h00;
 732 : data = 8'h00;
 733 : data = 8'h00;
 734 : data = 8'h00;
 735 : data = 8'h00;
 736 : data = 8'h00;
 737 : data = 8'h00;
 738 : data = 8'h00;
 739 : data = 8'h00;
 740 : data = 8'h00;
 741 : data = 8'h00;
 742 : data = 8'h00;
 743 : data = 8'h00;
 744 : data = 8'h00;
 745 : data = 8'h00;
 746 : data = 8'h00;
 747 : data = 8'h00;
 748 : data = 8'h00;
 749 : data = 8'h00;
 750 : data = 8'h00;
 751 : data = 8'h00;
 752 : data = 8'h00;
 753 : data = 8'h00;
 754 : data = 8'h00;
 755 : data = 8'h00;
 756 : data = 8'h00;
 757 : data = 8'h00;
 758 : data = 8'h00;
 759 : data = 8'h00;
 760 : data = 8'h00;
 761 : data = 8'h00;
 762 : data = 8'h00;
 763 : data = 8'h00;
 764 : data = 8'h00;
 765 : data = 8'h00;
 766 : data = 8'h00;
 767 : data = 8'h00;
 768 : data = 8'h00;
 769 : data = 8'h00;
 770 : data = 8'h00;
 771 : data = 8'h00;
 772 : data = 8'h00;
 773 : data = 8'h00;
 774 : data = 8'h00;
 775 : data = 8'h00;
 776 : data = 8'h00;
 777 : data = 8'h00;
 778 : data = 8'h00;
 779 : data = 8'h00;
 780 : data = 8'h00;
 781 : data = 8'h00;
 782 : data = 8'h00;
 783 : data = 8'h00;
 784 : data = 8'h00;
 785 : data = 8'h00;
 786 : data = 8'h00;
 787 : data = 8'h00;
 788 : data = 8'h00;
 789 : data = 8'h00;
 790 : data = 8'h00;
 791 : data = 8'h00;
 792 : data = 8'h00;
 793 : data = 8'h00;
 794 : data = 8'h00;
 795 : data = 8'h00;
 796 : data = 8'h00;
 797 : data = 8'h00;
 798 : data = 8'h00;
 799 : data = 8'h00;
 800 : data = 8'h00;
 801 : data = 8'h00;
 802 : data = 8'h00;
 803 : data = 8'h00;
 804 : data = 8'h00;
 805 : data = 8'h00;
 806 : data = 8'h00;
 807 : data = 8'h00;
 808 : data = 8'h00;
 809 : data = 8'h00;
 810 : data = 8'h00;
 811 : data = 8'h00;
 812 : data = 8'h00;
 813 : data = 8'h00;
 814 : data = 8'h00;
 815 : data = 8'h00;
 816 : data = 8'h00;
 817 : data = 8'h00;
 818 : data = 8'h00;
 819 : data = 8'h00;
 820 : data = 8'h00;
 821 : data = 8'h00;
 822 : data = 8'h00;
 823 : data = 8'h00;
 824 : data = 8'h00;
 825 : data = 8'h00;
 826 : data = 8'h00;
 827 : data = 8'h00;
 828 : data = 8'h00;
 829 : data = 8'h00;
 830 : data = 8'h00;
 831 : data = 8'h00;
 832 : data = 8'h00;
 833 : data = 8'h00;
 834 : data = 8'h00;
 835 : data = 8'h00;
 836 : data = 8'h00;
 837 : data = 8'h00;
 838 : data = 8'h00;
 839 : data = 8'h00;
 840 : data = 8'h00;
 841 : data = 8'h00;
 842 : data = 8'h00;
 843 : data = 8'h00;
 844 : data = 8'h00;
 845 : data = 8'h00;
 846 : data = 8'h00;
 847 : data = 8'h00;
 848 : data = 8'h00;
 849 : data = 8'h00;
 850 : data = 8'h00;
 851 : data = 8'h00;
 852 : data = 8'h00;
 853 : data = 8'h00;
 854 : data = 8'h00;
 855 : data = 8'h00;
 856 : data = 8'h00;
 857 : data = 8'h00;
 858 : data = 8'h00;
 859 : data = 8'h00;
 860 : data = 8'h00;
 861 : data = 8'h00;
 862 : data = 8'h00;
 863 : data = 8'h00;
 864 : data = 8'h00;
 865 : data = 8'h00;
 866 : data = 8'h00;
 867 : data = 8'h00;
 868 : data = 8'h00;
 869 : data = 8'h00;
 870 : data = 8'h00;
 871 : data = 8'h00;
 872 : data = 8'h00;
 873 : data = 8'h00;
 874 : data = 8'h00;
 875 : data = 8'h00;
 876 : data = 8'h00;
 877 : data = 8'h00;
 878 : data = 8'h00;
 879 : data = 8'h00;
 880 : data = 8'h00;
 881 : data = 8'h00;
 882 : data = 8'h00;
 883 : data = 8'h00;
 884 : data = 8'h00;
 885 : data = 8'h00;
 886 : data = 8'h00;
 887 : data = 8'h00;
 888 : data = 8'h00;
 889 : data = 8'h00;
 890 : data = 8'h00;
 891 : data = 8'h00;
 892 : data = 8'h00;
 893 : data = 8'h00;
 894 : data = 8'h00;
 895 : data = 8'h00;
 896 : data = 8'h00;
 897 : data = 8'h00;
 898 : data = 8'h00;
 899 : data = 8'h00;
 900 : data = 8'h00;
 901 : data = 8'h00;
 902 : data = 8'h00;
 903 : data = 8'h00;
 904 : data = 8'h00;
 905 : data = 8'h00;
 906 : data = 8'h00;
 907 : data = 8'h00;
 908 : data = 8'h00;
 909 : data = 8'h00;
 910 : data = 8'h00;
 911 : data = 8'h00;
 912 : data = 8'h00;
 913 : data = 8'h00;
 914 : data = 8'h00;
 915 : data = 8'h00;
 916 : data = 8'h00;
 917 : data = 8'h00;
 918 : data = 8'h00;
 919 : data = 8'h00;
 920 : data = 8'h00;
 921 : data = 8'h00;
 922 : data = 8'h00;
 923 : data = 8'h00;
 924 : data = 8'h00;
 925 : data = 8'h00;
 926 : data = 8'h00;
 927 : data = 8'h00;
 928 : data = 8'h00;
 929 : data = 8'h00;
 930 : data = 8'h00;
 931 : data = 8'h00;
 932 : data = 8'h00;
 933 : data = 8'h00;
 934 : data = 8'h00;
 935 : data = 8'h00;
 936 : data = 8'h00;
 937 : data = 8'h00;
 938 : data = 8'h00;
 939 : data = 8'h00;
 940 : data = 8'h00;
 941 : data = 8'h00;
 942 : data = 8'h00;
 943 : data = 8'h00;
 944 : data = 8'h00;
 945 : data = 8'h00;
 946 : data = 8'h00;
 947 : data = 8'h00;
 948 : data = 8'h00;
 949 : data = 8'h00;
 950 : data = 8'h00;
 951 : data = 8'h00;
 952 : data = 8'h00;
 953 : data = 8'h00;
 954 : data = 8'h00;
 955 : data = 8'h00;
 956 : data = 8'h00;
 957 : data = 8'h00;
 958 : data = 8'h00;
 959 : data = 8'h00;
 960 : data = 8'h00;
 961 : data = 8'h00;
 962 : data = 8'h00;
 963 : data = 8'h00;
 964 : data = 8'h00;
 965 : data = 8'h00;
 966 : data = 8'h00;
 967 : data = 8'h00;
 968 : data = 8'h00;
 969 : data = 8'h00;
 970 : data = 8'h00;
 971 : data = 8'h00;
 972 : data = 8'h00;
 973 : data = 8'h00;
 974 : data = 8'h00;
 975 : data = 8'h00;
 976 : data = 8'h00;
 977 : data = 8'h00;
 978 : data = 8'h00;
 979 : data = 8'h00;
 980 : data = 8'h00;
 981 : data = 8'h00;
 982 : data = 8'h00;
 983 : data = 8'h00;
 984 : data = 8'h00;
 985 : data = 8'h00;
 986 : data = 8'h00;
 987 : data = 8'h00;
 988 : data = 8'h00;
 989 : data = 8'h00;
 990 : data = 8'h00;
 991 : data = 8'h00;
 992 : data = 8'h00;
 993 : data = 8'h00;
 994 : data = 8'h00;
 995 : data = 8'h00;
 996 : data = 8'h00;
 997 : data = 8'h00;
 998 : data = 8'h00;
 999 : data = 8'h00;
 1000 : data = 8'h00;
 1001 : data = 8'h00;
 1002 : data = 8'h00;
 1003 : data = 8'h00;
 1004 : data = 8'h00;
 1005 : data = 8'h00;
 1006 : data = 8'h00;
 1007 : data = 8'h00;
 1008 : data = 8'h00;
 1009 : data = 8'h00;
 1010 : data = 8'h00;
 1011 : data = 8'h00;
 1012 : data = 8'h00;
 1013 : data = 8'h00;
 1014 : data = 8'h00;
 1015 : data = 8'h00;
 1016 : data = 8'h00;
 1017 : data = 8'h00;
 1018 : data = 8'h00;
 1019 : data = 8'h00;
 1020 : data = 8'h00;
 1021 : data = 8'h00;
 1022 : data = 8'h00;
 1023 : data = 8'h00;
 1024 : data = 8'h00;
 1025 : data = 8'h00;
 1026 : data = 8'h00;
 1027 : data = 8'h00;
 1028 : data = 8'h00;
 1029 : data = 8'h00;
 1030 : data = 8'h00;
 1031 : data = 8'h00;
 1032 : data = 8'h00;
 1033 : data = 8'h00;
 1034 : data = 8'h00;
 1035 : data = 8'h00;
 1036 : data = 8'h00;
 1037 : data = 8'h00;
 1038 : data = 8'h00;
 1039 : data = 8'h00;
 1040 : data = 8'h00;
 1041 : data = 8'h00;
 1042 : data = 8'h00;
 1043 : data = 8'h00;
 1044 : data = 8'h00;
 1045 : data = 8'h00;
 1046 : data = 8'h00;
 1047 : data = 8'h00;
 1048 : data = 8'h00;
 1049 : data = 8'h00;
 1050 : data = 8'h00;
 1051 : data = 8'h00;
 1052 : data = 8'h00;
 1053 : data = 8'h00;
 1054 : data = 8'h00;
 1055 : data = 8'h00;
 1056 : data = 8'h00;
 1057 : data = 8'h00;
 1058 : data = 8'h00;
 1059 : data = 8'h00;
 1060 : data = 8'h00;
 1061 : data = 8'h00;
 1062 : data = 8'h00;
 1063 : data = 8'h00;
 1064 : data = 8'h00;
 1065 : data = 8'h00;
 1066 : data = 8'h00;
 1067 : data = 8'h00;
 1068 : data = 8'h00;
 1069 : data = 8'h00;
 1070 : data = 8'h00;
 1071 : data = 8'h00;
 1072 : data = 8'h00;
 1073 : data = 8'h00;
 1074 : data = 8'h00;
 1075 : data = 8'h00;
 1076 : data = 8'h00;
 1077 : data = 8'h00;
 1078 : data = 8'h00;
 1079 : data = 8'h00;
 1080 : data = 8'h00;
 1081 : data = 8'h00;
 1082 : data = 8'h00;
 1083 : data = 8'h00;
 1084 : data = 8'h00;
 1085 : data = 8'h00;
 1086 : data = 8'h00;
 1087 : data = 8'h00;
 1088 : data = 8'h00;
 1089 : data = 8'h00;
 1090 : data = 8'h00;
 1091 : data = 8'h00;
 1092 : data = 8'h00;
 1093 : data = 8'h00;
 1094 : data = 8'h00;
 1095 : data = 8'h00;
 1096 : data = 8'h00;
 1097 : data = 8'h00;
 1098 : data = 8'h00;
 1099 : data = 8'h00;
 1100 : data = 8'h00;
 1101 : data = 8'h00;
 1102 : data = 8'h00;
 1103 : data = 8'h00;
 1104 : data = 8'h00;
 1105 : data = 8'h00;
 1106 : data = 8'h00;
 1107 : data = 8'h00;
 1108 : data = 8'h00;
 1109 : data = 8'h00;
 1110 : data = 8'h00;
 1111 : data = 8'h00;
 1112 : data = 8'h00;
 1113 : data = 8'h00;
 1114 : data = 8'h00;
 1115 : data = 8'h00;
 1116 : data = 8'h00;
 1117 : data = 8'h00;
 1118 : data = 8'h00;
 1119 : data = 8'h00;
 1120 : data = 8'h00;
 1121 : data = 8'h00;
 1122 : data = 8'h00;
 1123 : data = 8'h00;
 1124 : data = 8'h00;
 1125 : data = 8'h00;
 1126 : data = 8'h00;
 1127 : data = 8'h00;
 1128 : data = 8'h00;
 1129 : data = 8'h00;
 1130 : data = 8'h00;
 1131 : data = 8'h00;
 1132 : data = 8'h00;
 1133 : data = 8'h00;
 1134 : data = 8'h00;
 1135 : data = 8'h00;
 1136 : data = 8'h00;
 1137 : data = 8'h00;
 1138 : data = 8'h00;
 1139 : data = 8'h00;
 1140 : data = 8'h00;
 1141 : data = 8'h00;
 1142 : data = 8'h00;
 1143 : data = 8'h00;
 1144 : data = 8'h00;
 1145 : data = 8'h00;
 1146 : data = 8'h00;
 1147 : data = 8'h00;
 1148 : data = 8'h00;
 1149 : data = 8'h00;
 1150 : data = 8'h00;
 1151 : data = 8'h00;
 1152 : data = 8'h00;
 1153 : data = 8'h00;
 1154 : data = 8'h00;
 1155 : data = 8'h00;
 1156 : data = 8'h00;
 1157 : data = 8'h00;
 1158 : data = 8'h00;
 1159 : data = 8'h00;
 1160 : data = 8'h00;
 1161 : data = 8'h00;
 1162 : data = 8'h00;
 1163 : data = 8'h00;
 1164 : data = 8'h00;
 1165 : data = 8'h00;
 1166 : data = 8'h00;
 1167 : data = 8'h00;
 1168 : data = 8'h00;
 1169 : data = 8'h00;
 1170 : data = 8'h00;
 1171 : data = 8'h00;
 1172 : data = 8'h00;
 1173 : data = 8'h00;
 1174 : data = 8'h00;
 1175 : data = 8'h00;
 1176 : data = 8'h00;
 1177 : data = 8'h00;
 1178 : data = 8'h00;
 1179 : data = 8'h00;
 1180 : data = 8'h00;
 1181 : data = 8'h00;
 1182 : data = 8'h00;
 1183 : data = 8'h00;
 1184 : data = 8'h00;
 1185 : data = 8'h00;
 1186 : data = 8'h00;
 1187 : data = 8'h00;
 1188 : data = 8'h00;
 1189 : data = 8'h00;
 1190 : data = 8'h00;
 1191 : data = 8'h00;
 1192 : data = 8'h00;
 1193 : data = 8'h00;
 1194 : data = 8'h00;
 1195 : data = 8'h00;
 1196 : data = 8'h00;
 1197 : data = 8'h00;
 1198 : data = 8'h00;
 1199 : data = 8'h00;
 1200 : data = 8'h00;
 1201 : data = 8'h00;
 1202 : data = 8'h00;
 1203 : data = 8'h00;
 1204 : data = 8'h00;
 1205 : data = 8'h00;
 1206 : data = 8'h00;
 1207 : data = 8'h00;
 1208 : data = 8'h00;
 1209 : data = 8'h00;
 1210 : data = 8'h00;
 1211 : data = 8'h00;
 1212 : data = 8'h00;
 1213 : data = 8'h00;
 1214 : data = 8'h00;
 1215 : data = 8'h00;
 1216 : data = 8'h00;
 1217 : data = 8'h00;
 1218 : data = 8'h00;
 1219 : data = 8'h00;
 1220 : data = 8'h00;
 1221 : data = 8'h00;
 1222 : data = 8'h00;
 1223 : data = 8'h00;
 1224 : data = 8'h00;
 1225 : data = 8'h00;
 1226 : data = 8'h00;
 1227 : data = 8'h00;
 1228 : data = 8'h00;
 1229 : data = 8'h00;
 1230 : data = 8'h00;
 1231 : data = 8'h00;
 1232 : data = 8'h00;
 1233 : data = 8'h00;
 1234 : data = 8'h00;
 1235 : data = 8'h00;
 1236 : data = 8'h00;
 1237 : data = 8'h00;
 1238 : data = 8'h00;
 1239 : data = 8'h00;
 1240 : data = 8'h00;
 1241 : data = 8'h00;
 1242 : data = 8'h00;
 1243 : data = 8'h00;
 1244 : data = 8'h00;
 1245 : data = 8'h00;
 1246 : data = 8'h00;
 1247 : data = 8'h00;
 1248 : data = 8'h00;
 1249 : data = 8'h00;
 1250 : data = 8'h00;
 1251 : data = 8'h00;
 1252 : data = 8'h00;
 1253 : data = 8'h00;
 1254 : data = 8'h00;
 1255 : data = 8'h00;
 1256 : data = 8'h00;
 1257 : data = 8'h00;
 1258 : data = 8'h00;
 1259 : data = 8'h00;
 1260 : data = 8'h00;
 1261 : data = 8'h00;
 1262 : data = 8'h00;
 1263 : data = 8'h00;
 1264 : data = 8'h00;
 1265 : data = 8'h00;
 1266 : data = 8'h00;
 1267 : data = 8'h00;
 1268 : data = 8'h00;
 1269 : data = 8'h00;
 1270 : data = 8'h00;
 1271 : data = 8'h00;
 1272 : data = 8'h00;
 1273 : data = 8'h00;
 1274 : data = 8'h00;
 1275 : data = 8'h00;
 1276 : data = 8'h00;
 1277 : data = 8'h00;
 1278 : data = 8'h00;
 1279 : data = 8'h00;
 1280 : data = 8'h00;
 1281 : data = 8'h00;
 1282 : data = 8'h00;
 1283 : data = 8'h00;
 1284 : data = 8'h00;
 1285 : data = 8'h00;
 1286 : data = 8'h00;
 1287 : data = 8'h00;
 1288 : data = 8'h00;
 1289 : data = 8'h00;
 1290 : data = 8'h00;
 1291 : data = 8'h00;
 1292 : data = 8'h00;
 1293 : data = 8'h00;
 1294 : data = 8'h00;
 1295 : data = 8'h00;
 1296 : data = 8'h00;
 1297 : data = 8'h00;
 1298 : data = 8'h00;
 1299 : data = 8'h00;
 1300 : data = 8'h00;
 1301 : data = 8'h00;
 1302 : data = 8'h00;
 1303 : data = 8'h00;
 1304 : data = 8'h00;
 1305 : data = 8'h00;
 1306 : data = 8'h00;
 1307 : data = 8'h00;
 1308 : data = 8'h00;
 1309 : data = 8'h00;
 1310 : data = 8'h00;
 1311 : data = 8'h00;
 1312 : data = 8'h00;
 1313 : data = 8'h00;
 1314 : data = 8'h00;
 1315 : data = 8'h00;
 1316 : data = 8'h00;
 1317 : data = 8'h00;
 1318 : data = 8'h00;
 1319 : data = 8'h00;
 1320 : data = 8'h00;
 1321 : data = 8'h00;
 1322 : data = 8'h00;
 1323 : data = 8'h00;
 1324 : data = 8'h00;
 1325 : data = 8'h00;
 1326 : data = 8'h00;
 1327 : data = 8'h00;
 1328 : data = 8'h00;
 1329 : data = 8'h00;
 1330 : data = 8'h00;
 1331 : data = 8'h00;
 1332 : data = 8'h00;
 1333 : data = 8'h00;
 1334 : data = 8'h00;
 1335 : data = 8'h00;
 1336 : data = 8'h00;
 1337 : data = 8'h00;
 1338 : data = 8'h00;
 1339 : data = 8'h00;
 1340 : data = 8'h00;
 1341 : data = 8'h00;
 1342 : data = 8'h00;
 1343 : data = 8'h00;
 1344 : data = 8'h00;
 1345 : data = 8'h00;
 1346 : data = 8'h00;
 1347 : data = 8'h00;
 1348 : data = 8'h00;
 1349 : data = 8'h00;
 1350 : data = 8'h00;
 1351 : data = 8'h00;
 1352 : data = 8'h00;
 1353 : data = 8'h00;
 1354 : data = 8'h00;
 1355 : data = 8'h00;
 1356 : data = 8'h00;
 1357 : data = 8'h00;
 1358 : data = 8'h00;
 1359 : data = 8'h00;
 1360 : data = 8'h00;
 1361 : data = 8'h00;
 1362 : data = 8'h00;
 1363 : data = 8'h00;
 1364 : data = 8'h00;
 1365 : data = 8'h00;
 1366 : data = 8'h00;
 1367 : data = 8'h00;
 1368 : data = 8'h00;
 1369 : data = 8'h00;
 1370 : data = 8'h00;
 1371 : data = 8'h00;
 1372 : data = 8'h00;
 1373 : data = 8'h00;
 1374 : data = 8'h00;
 1375 : data = 8'h00;
 1376 : data = 8'h00;
 1377 : data = 8'h00;
 1378 : data = 8'h00;
 1379 : data = 8'h00;
 1380 : data = 8'h00;
 1381 : data = 8'h00;
 1382 : data = 8'h00;
 1383 : data = 8'h00;
 1384 : data = 8'h00;
 1385 : data = 8'h00;
 1386 : data = 8'h00;
 1387 : data = 8'h00;
 1388 : data = 8'h00;
 1389 : data = 8'h00;
 1390 : data = 8'h00;
 1391 : data = 8'h00;
 1392 : data = 8'h00;
 1393 : data = 8'h00;
 1394 : data = 8'h00;
 1395 : data = 8'h00;
 1396 : data = 8'h00;
 1397 : data = 8'h00;
 1398 : data = 8'h00;
 1399 : data = 8'h00;
 1400 : data = 8'h00;
 1401 : data = 8'h00;
 1402 : data = 8'h00;
 1403 : data = 8'h00;
 1404 : data = 8'h00;
 1405 : data = 8'h00;
 1406 : data = 8'h00;
 1407 : data = 8'h00;
 1408 : data = 8'h00;
 1409 : data = 8'h00;
 1410 : data = 8'h00;
 1411 : data = 8'h00;
 1412 : data = 8'h00;
 1413 : data = 8'h00;
 1414 : data = 8'h00;
 1415 : data = 8'h00;
 1416 : data = 8'h00;
 1417 : data = 8'h00;
 1418 : data = 8'h00;
 1419 : data = 8'h00;
 1420 : data = 8'h00;
 1421 : data = 8'h00;
 1422 : data = 8'h00;
 1423 : data = 8'h00;
 1424 : data = 8'h00;
 1425 : data = 8'h00;
 1426 : data = 8'h00;
 1427 : data = 8'h00;
 1428 : data = 8'h00;
 1429 : data = 8'h00;
 1430 : data = 8'h00;
 1431 : data = 8'h00;
 1432 : data = 8'h00;
 1433 : data = 8'h00;
 1434 : data = 8'h00;
 1435 : data = 8'h00;
 1436 : data = 8'h00;
 1437 : data = 8'h00;
 1438 : data = 8'h00;
 1439 : data = 8'h00;
 1440 : data = 8'h00;
 1441 : data = 8'h00;
 1442 : data = 8'h00;
 1443 : data = 8'h00;
 1444 : data = 8'h00;
 1445 : data = 8'h00;
 1446 : data = 8'h00;
 1447 : data = 8'h00;
 1448 : data = 8'h00;
 1449 : data = 8'h00;
 1450 : data = 8'h00;
 1451 : data = 8'h00;
 1452 : data = 8'h00;
 1453 : data = 8'h00;
 1454 : data = 8'h00;
 1455 : data = 8'h00;
 1456 : data = 8'h00;
 1457 : data = 8'h00;
 1458 : data = 8'h00;
 1459 : data = 8'h00;
 1460 : data = 8'h00;
 1461 : data = 8'h00;
 1462 : data = 8'h00;
 1463 : data = 8'h00;
 1464 : data = 8'h00;
 1465 : data = 8'h00;
 1466 : data = 8'h00;
 1467 : data = 8'h00;
 1468 : data = 8'h00;
 1469 : data = 8'h00;
 1470 : data = 8'h00;
 1471 : data = 8'h00;
 1472 : data = 8'h00;
 1473 : data = 8'h00;
 1474 : data = 8'h00;
 1475 : data = 8'h00;
 1476 : data = 8'h00;
 1477 : data = 8'h00;
 1478 : data = 8'h00;
 1479 : data = 8'h00;
 1480 : data = 8'h00;
 1481 : data = 8'h00;
 1482 : data = 8'h00;
 1483 : data = 8'h00;
 1484 : data = 8'h00;
 1485 : data = 8'h00;
 1486 : data = 8'h00;
 1487 : data = 8'h00;
 1488 : data = 8'h00;
 1489 : data = 8'h00;
 1490 : data = 8'h00;
 1491 : data = 8'h00;
 1492 : data = 8'h00;
 1493 : data = 8'h00;
 1494 : data = 8'h00;
 1495 : data = 8'h00;
 1496 : data = 8'h00;
 1497 : data = 8'h00;
 1498 : data = 8'h00;
 1499 : data = 8'h00;
 1500 : data = 8'h00;
 1501 : data = 8'h00;
 1502 : data = 8'h00;
 1503 : data = 8'h00;
 1504 : data = 8'h00;
 1505 : data = 8'h00;
 1506 : data = 8'h00;
 1507 : data = 8'h00;
 1508 : data = 8'h00;
 1509 : data = 8'h00;
 1510 : data = 8'h00;
 1511 : data = 8'h00;
 1512 : data = 8'h00;
 1513 : data = 8'h00;
 1514 : data = 8'h00;
 1515 : data = 8'h00;
 1516 : data = 8'h00;
 1517 : data = 8'h00;
 1518 : data = 8'h00;
 1519 : data = 8'h00;
 1520 : data = 8'h00;
 1521 : data = 8'h00;
 1522 : data = 8'h00;
 1523 : data = 8'h00;
 1524 : data = 8'h00;
 1525 : data = 8'h00;
 1526 : data = 8'h00;
 1527 : data = 8'h00;
 1528 : data = 8'h00;
 1529 : data = 8'h00;
 1530 : data = 8'h00;
 1531 : data = 8'h00;
 1532 : data = 8'h00;
 1533 : data = 8'h00;
 1534 : data = 8'h00;
 1535 : data = 8'h00;
 1536 : data = 8'h00;
 1537 : data = 8'h00;
 1538 : data = 8'h00;
 1539 : data = 8'h00;
 1540 : data = 8'h00;
 1541 : data = 8'h00;
 1542 : data = 8'h00;
 1543 : data = 8'h00;
 1544 : data = 8'h00;
 1545 : data = 8'h00;
 1546 : data = 8'h00;
 1547 : data = 8'h00;
 1548 : data = 8'h00;
 1549 : data = 8'h00;
 1550 : data = 8'h00;
 1551 : data = 8'h00;
 1552 : data = 8'h00;
 1553 : data = 8'h00;
 1554 : data = 8'h00;
 1555 : data = 8'h00;
 1556 : data = 8'h00;
 1557 : data = 8'h00;
 1558 : data = 8'h00;
 1559 : data = 8'h00;
 1560 : data = 8'h00;
 1561 : data = 8'h00;
 1562 : data = 8'h00;
 1563 : data = 8'h00;
 1564 : data = 8'h00;
 1565 : data = 8'h00;
 1566 : data = 8'h00;
 1567 : data = 8'h00;
 1568 : data = 8'h00;
 1569 : data = 8'h00;
 1570 : data = 8'h00;
 1571 : data = 8'h00;
 1572 : data = 8'h00;
 1573 : data = 8'h00;
 1574 : data = 8'h00;
 1575 : data = 8'h00;
 1576 : data = 8'h00;
 1577 : data = 8'h00;
 1578 : data = 8'h00;
 1579 : data = 8'h00;
 1580 : data = 8'h00;
 1581 : data = 8'h00;
 1582 : data = 8'h00;
 1583 : data = 8'h00;
 1584 : data = 8'h00;
 1585 : data = 8'h00;
 1586 : data = 8'h00;
 1587 : data = 8'h00;
 1588 : data = 8'h00;
 1589 : data = 8'h00;
 1590 : data = 8'h00;
 1591 : data = 8'h00;
 1592 : data = 8'h00;
 1593 : data = 8'h00;
 1594 : data = 8'h00;
 1595 : data = 8'h00;
 1596 : data = 8'h00;
 1597 : data = 8'h00;
 1598 : data = 8'h00;
 1599 : data = 8'h00;
 1600 : data = 8'h00;
 1601 : data = 8'h00;
 1602 : data = 8'h00;
 1603 : data = 8'h00;
 1604 : data = 8'h00;
 1605 : data = 8'h00;
 1606 : data = 8'h00;
 1607 : data = 8'h00;
 1608 : data = 8'h00;
 1609 : data = 8'h00;
 1610 : data = 8'h00;
 1611 : data = 8'h00;
 1612 : data = 8'h00;
 1613 : data = 8'h00;
 1614 : data = 8'h00;
 1615 : data = 8'h00;
 1616 : data = 8'h00;
 1617 : data = 8'h00;
 1618 : data = 8'h00;
 1619 : data = 8'h00;
 1620 : data = 8'h00;
 1621 : data = 8'h00;
 1622 : data = 8'h00;
 1623 : data = 8'h00;
 1624 : data = 8'h00;
 1625 : data = 8'h00;
 1626 : data = 8'h00;
 1627 : data = 8'h00;
 1628 : data = 8'h00;
 1629 : data = 8'h00;
 1630 : data = 8'h00;
 1631 : data = 8'h00;
 1632 : data = 8'h00;
 1633 : data = 8'h00;
 1634 : data = 8'h00;
 1635 : data = 8'h00;
 1636 : data = 8'h00;
 1637 : data = 8'h00;
 1638 : data = 8'h00;
 1639 : data = 8'h00;
 1640 : data = 8'h00;
 1641 : data = 8'h00;
 1642 : data = 8'h00;
 1643 : data = 8'h00;
 1644 : data = 8'h00;
 1645 : data = 8'h00;
 1646 : data = 8'h00;
 1647 : data = 8'h00;
 1648 : data = 8'h00;
 1649 : data = 8'h00;
 1650 : data = 8'h00;
 1651 : data = 8'h00;
 1652 : data = 8'h00;
 1653 : data = 8'h00;
 1654 : data = 8'h00;
 1655 : data = 8'h00;
 1656 : data = 8'h00;
 1657 : data = 8'h00;
 1658 : data = 8'h00;
 1659 : data = 8'h00;
 1660 : data = 8'h00;
 1661 : data = 8'h00;
 1662 : data = 8'h00;
 1663 : data = 8'h00;
 1664 : data = 8'h00;
 1665 : data = 8'h00;
 1666 : data = 8'h00;
 1667 : data = 8'h00;
 1668 : data = 8'h00;
 1669 : data = 8'h00;
 1670 : data = 8'h00;
 1671 : data = 8'h00;
 1672 : data = 8'h00;
 1673 : data = 8'h00;
 1674 : data = 8'h00;
 1675 : data = 8'h00;
 1676 : data = 8'h00;
 1677 : data = 8'h00;
 1678 : data = 8'h00;
 1679 : data = 8'h00;
 1680 : data = 8'h00;
 1681 : data = 8'h00;
 1682 : data = 8'h00;
 1683 : data = 8'h00;
 1684 : data = 8'h00;
 1685 : data = 8'h00;
 1686 : data = 8'h00;
 1687 : data = 8'h00;
 1688 : data = 8'h00;
 1689 : data = 8'h00;
 1690 : data = 8'h00;
 1691 : data = 8'h00;
 1692 : data = 8'h00;
 1693 : data = 8'h00;
 1694 : data = 8'h00;
 1695 : data = 8'h00;
 1696 : data = 8'h00;
 1697 : data = 8'h00;
 1698 : data = 8'h00;
 1699 : data = 8'h00;
 1700 : data = 8'h00;
 1701 : data = 8'h00;
 1702 : data = 8'h00;
 1703 : data = 8'h00;
 1704 : data = 8'h00;
 1705 : data = 8'h00;
 1706 : data = 8'h00;
 1707 : data = 8'h00;
 1708 : data = 8'h00;
 1709 : data = 8'h00;
 1710 : data = 8'h00;
 1711 : data = 8'h00;
 1712 : data = 8'h00;
 1713 : data = 8'h00;
 1714 : data = 8'h00;
 1715 : data = 8'h00;
 1716 : data = 8'h00;
 1717 : data = 8'h00;
 1718 : data = 8'h00;
 1719 : data = 8'h00;
 1720 : data = 8'h00;
 1721 : data = 8'h00;
 1722 : data = 8'h00;
 1723 : data = 8'h00;
 1724 : data = 8'h00;
 1725 : data = 8'h00;
 1726 : data = 8'h00;
 1727 : data = 8'h00;
 1728 : data = 8'h00;
 1729 : data = 8'h00;
 1730 : data = 8'h00;
 1731 : data = 8'h00;
 1732 : data = 8'h00;
 1733 : data = 8'h00;
 1734 : data = 8'h00;
 1735 : data = 8'h00;
 1736 : data = 8'h00;
 1737 : data = 8'h00;
 1738 : data = 8'h00;
 1739 : data = 8'h00;
 1740 : data = 8'h00;
 1741 : data = 8'h00;
 1742 : data = 8'h00;
 1743 : data = 8'h00;
 1744 : data = 8'h00;
 1745 : data = 8'h00;
 1746 : data = 8'h00;
 1747 : data = 8'h00;
 1748 : data = 8'h00;
 1749 : data = 8'h00;
 1750 : data = 8'h00;
 1751 : data = 8'h00;
 1752 : data = 8'h00;
 1753 : data = 8'h00;
 1754 : data = 8'h00;
 1755 : data = 8'h00;
 1756 : data = 8'h00;
 1757 : data = 8'h00;
 1758 : data = 8'h00;
 1759 : data = 8'h00;
 1760 : data = 8'h00;
 1761 : data = 8'h00;
 1762 : data = 8'h00;
 1763 : data = 8'h00;
 1764 : data = 8'h00;
 1765 : data = 8'h00;
 1766 : data = 8'h00;
 1767 : data = 8'h00;
 1768 : data = 8'h00;
 1769 : data = 8'h00;
 1770 : data = 8'h00;
 1771 : data = 8'h00;
 1772 : data = 8'h00;
 1773 : data = 8'h00;
 1774 : data = 8'h00;
 1775 : data = 8'h00;
 1776 : data = 8'h00;
 1777 : data = 8'h00;
 1778 : data = 8'h00;
 1779 : data = 8'h00;
 1780 : data = 8'h00;
 1781 : data = 8'h00;
 1782 : data = 8'h00;
 1783 : data = 8'h00;
 1784 : data = 8'h00;
 1785 : data = 8'h00;
 1786 : data = 8'h00;
 1787 : data = 8'h00;
 1788 : data = 8'h00;
 1789 : data = 8'h00;
 1790 : data = 8'h00;
 1791 : data = 8'h00;
 1792 : data = 8'h00;
 1793 : data = 8'h00;
 1794 : data = 8'h00;
 1795 : data = 8'h00;
 1796 : data = 8'h00;
 1797 : data = 8'h00;
 1798 : data = 8'h00;
 1799 : data = 8'h00;
 1800 : data = 8'h00;
 1801 : data = 8'h00;
 1802 : data = 8'h00;
 1803 : data = 8'h00;
 1804 : data = 8'h00;
 1805 : data = 8'h00;
 1806 : data = 8'h00;
 1807 : data = 8'h00;
 1808 : data = 8'h00;
 1809 : data = 8'h00;
 1810 : data = 8'h00;
 1811 : data = 8'h00;
 1812 : data = 8'h00;
 1813 : data = 8'h00;
 1814 : data = 8'h00;
 1815 : data = 8'h00;
 1816 : data = 8'h00;
 1817 : data = 8'h00;
 1818 : data = 8'h00;
 1819 : data = 8'h00;
 1820 : data = 8'h00;
 1821 : data = 8'h00;
 1822 : data = 8'h00;
 1823 : data = 8'h00;
 1824 : data = 8'h00;
 1825 : data = 8'h00;
 1826 : data = 8'h00;
 1827 : data = 8'h00;
 1828 : data = 8'h00;
 1829 : data = 8'h00;
 1830 : data = 8'h00;
 1831 : data = 8'h00;
 1832 : data = 8'h00;
 1833 : data = 8'h00;
 1834 : data = 8'h00;
 1835 : data = 8'h00;
 1836 : data = 8'h00;
 1837 : data = 8'h00;
 1838 : data = 8'h00;
 1839 : data = 8'h00;
 1840 : data = 8'h00;
 1841 : data = 8'h00;
 1842 : data = 8'h00;
 1843 : data = 8'h00;
 1844 : data = 8'h00;
 1845 : data = 8'h00;
 1846 : data = 8'h00;
 1847 : data = 8'h00;
 1848 : data = 8'h00;
 1849 : data = 8'h00;
 1850 : data = 8'h00;
 1851 : data = 8'h00;
 1852 : data = 8'h00;
 1853 : data = 8'h00;
 1854 : data = 8'h00;
 1855 : data = 8'h00;
 1856 : data = 8'h00;
 1857 : data = 8'h00;
 1858 : data = 8'h00;
 1859 : data = 8'h00;
 1860 : data = 8'h00;
 1861 : data = 8'h00;
 1862 : data = 8'h00;
 1863 : data = 8'h00;
 1864 : data = 8'h00;
 1865 : data = 8'h00;
 1866 : data = 8'h00;
 1867 : data = 8'h00;
 1868 : data = 8'h00;
 1869 : data = 8'h00;
 1870 : data = 8'h00;
 1871 : data = 8'h00;
 1872 : data = 8'h00;
 1873 : data = 8'h00;
 1874 : data = 8'h00;
 1875 : data = 8'h00;
 1876 : data = 8'h00;
 1877 : data = 8'h00;
 1878 : data = 8'h00;
 1879 : data = 8'h00;
 1880 : data = 8'h00;
 1881 : data = 8'h00;
 1882 : data = 8'h00;
 1883 : data = 8'h00;
 1884 : data = 8'h00;
 1885 : data = 8'h00;
 1886 : data = 8'h00;
 1887 : data = 8'h00;
 1888 : data = 8'h00;
 1889 : data = 8'h00;
 1890 : data = 8'h00;
 1891 : data = 8'h00;
 1892 : data = 8'h00;
 1893 : data = 8'h00;
 1894 : data = 8'h00;
 1895 : data = 8'h00;
 1896 : data = 8'h00;
 1897 : data = 8'h00;
 1898 : data = 8'h00;
 1899 : data = 8'h00;
 1900 : data = 8'h00;
 1901 : data = 8'h00;
 1902 : data = 8'h00;
 1903 : data = 8'h00;
 1904 : data = 8'h00;
 1905 : data = 8'h00;
 1906 : data = 8'h00;
 1907 : data = 8'h00;
 1908 : data = 8'h00;
 1909 : data = 8'h00;
 1910 : data = 8'h00;
 1911 : data = 8'h00;
 1912 : data = 8'h00;
 1913 : data = 8'h00;
 1914 : data = 8'h00;
 1915 : data = 8'h00;
 1916 : data = 8'h00;
 1917 : data = 8'h00;
 1918 : data = 8'h00;
 1919 : data = 8'h00;
 1920 : data = 8'h00;
 1921 : data = 8'h00;
 1922 : data = 8'h00;
 1923 : data = 8'h00;
 1924 : data = 8'h00;
 1925 : data = 8'h00;
 1926 : data = 8'h00;
 1927 : data = 8'h00;
 1928 : data = 8'h00;
 1929 : data = 8'h00;
 1930 : data = 8'h00;
 1931 : data = 8'h00;
 1932 : data = 8'h00;
 1933 : data = 8'h00;
 1934 : data = 8'h00;
 1935 : data = 8'h00;
 1936 : data = 8'h00;
 1937 : data = 8'h00;
 1938 : data = 8'h00;
 1939 : data = 8'h00;
 1940 : data = 8'h00;
 1941 : data = 8'h00;
 1942 : data = 8'h00;
 1943 : data = 8'h00;
 1944 : data = 8'h00;
 1945 : data = 8'h00;
 1946 : data = 8'h00;
 1947 : data = 8'h00;
 1948 : data = 8'h00;
 1949 : data = 8'h00;
 1950 : data = 8'h00;
 1951 : data = 8'h00;
 1952 : data = 8'h00;
 1953 : data = 8'h00;
 1954 : data = 8'h00;
 1955 : data = 8'h00;
 1956 : data = 8'h00;
 1957 : data = 8'h00;
 1958 : data = 8'h00;
 1959 : data = 8'h00;
 1960 : data = 8'h00;
 1961 : data = 8'h00;
 1962 : data = 8'h00;
 1963 : data = 8'h00;
 1964 : data = 8'h00;
 1965 : data = 8'h00;
 1966 : data = 8'h00;
 1967 : data = 8'h00;
 1968 : data = 8'h00;
 1969 : data = 8'h00;
 1970 : data = 8'h00;
 1971 : data = 8'h00;
 1972 : data = 8'h00;
 1973 : data = 8'h00;
 1974 : data = 8'h00;
 1975 : data = 8'h00;
 1976 : data = 8'h00;
 1977 : data = 8'h00;
 1978 : data = 8'h00;
 1979 : data = 8'h00;
 1980 : data = 8'h00;
 1981 : data = 8'h00;
 1982 : data = 8'h00;
 1983 : data = 8'h00;
 1984 : data = 8'h00;
 1985 : data = 8'h00;
 1986 : data = 8'h00;
 1987 : data = 8'h00;
 1988 : data = 8'h00;
 1989 : data = 8'h00;
 1990 : data = 8'h00;
 1991 : data = 8'h00;
 1992 : data = 8'h00;
 1993 : data = 8'h00;
 1994 : data = 8'h00;
 1995 : data = 8'h00;
 1996 : data = 8'h00;
 1997 : data = 8'h00;
 1998 : data = 8'h00;
 1999 : data = 8'h00;
 2000 : data = 8'h00;
 2001 : data = 8'h00;
 2002 : data = 8'h00;
 2003 : data = 8'h00;
 2004 : data = 8'h00;
 2005 : data = 8'h00;
 2006 : data = 8'h00;
 2007 : data = 8'h00;
 2008 : data = 8'h00;
 2009 : data = 8'h00;
 2010 : data = 8'h00;
 2011 : data = 8'h00;
 2012 : data = 8'h00;
 2013 : data = 8'h00;
 2014 : data = 8'h00;
 2015 : data = 8'h00;
 2016 : data = 8'h00;
 2017 : data = 8'h00;
 2018 : data = 8'h00;
 2019 : data = 8'h00;
 2020 : data = 8'h00;
 2021 : data = 8'h00;
 2022 : data = 8'h00;
 2023 : data = 8'h00;
 2024 : data = 8'h00;
 2025 : data = 8'h00;
 2026 : data = 8'h00;
 2027 : data = 8'h00;
 2028 : data = 8'h00;
 2029 : data = 8'h00;
 2030 : data = 8'h00;
 2031 : data = 8'h00;
 2032 : data = 8'h00;
 2033 : data = 8'h00;
 2034 : data = 8'h00;
 2035 : data = 8'h00;
 2036 : data = 8'h00;
 2037 : data = 8'h00;
 2038 : data = 8'h00;
 2039 : data = 8'h00;
 2040 : data = 8'h00;
 2041 : data = 8'h00;
 2042 : data = 8'h00;
 2043 : data = 8'h00;
 2044 : data = 8'h00;
 2045 : data = 8'h00;
 2046 : data = 8'h00;
 2047 : data = 8'h00;
 2048 : data = 8'h00;
 2049 : data = 8'h00;
 2050 : data = 8'h00;
 2051 : data = 8'h00;
 2052 : data = 8'h00;
 2053 : data = 8'h00;
 2054 : data = 8'h00;
 2055 : data = 8'h00;
 2056 : data = 8'h00;
 2057 : data = 8'h00;
 2058 : data = 8'h00;
 2059 : data = 8'h00;
 2060 : data = 8'h00;
 2061 : data = 8'h00;
 2062 : data = 8'h00;
 2063 : data = 8'h00;
 2064 : data = 8'h00;
 2065 : data = 8'h00;
 2066 : data = 8'h00;
 2067 : data = 8'h00;
 2068 : data = 8'h00;
 2069 : data = 8'h00;
 2070 : data = 8'h00;
 2071 : data = 8'h00;
 2072 : data = 8'h00;
 2073 : data = 8'h00;
 2074 : data = 8'h00;
 2075 : data = 8'h00;
 2076 : data = 8'h00;
 2077 : data = 8'h00;
 2078 : data = 8'h00;
 2079 : data = 8'h00;
 2080 : data = 8'h00;
 2081 : data = 8'h00;
 2082 : data = 8'h00;
 2083 : data = 8'h00;
 2084 : data = 8'h00;
 2085 : data = 8'h00;
 2086 : data = 8'h00;
 2087 : data = 8'h00;
 2088 : data = 8'h00;
 2089 : data = 8'h00;
 2090 : data = 8'h00;
 2091 : data = 8'h00;
 2092 : data = 8'h00;
 2093 : data = 8'h00;
 2094 : data = 8'h00;
 2095 : data = 8'h00;
 2096 : data = 8'h00;
 2097 : data = 8'h00;
 2098 : data = 8'h00;
 2099 : data = 8'h00;
 2100 : data = 8'h00;
 2101 : data = 8'h00;
 2102 : data = 8'h00;
 2103 : data = 8'h00;
 2104 : data = 8'h00;
 2105 : data = 8'h00;
 2106 : data = 8'h00;
 2107 : data = 8'h00;
 2108 : data = 8'h00;
 2109 : data = 8'h00;
 2110 : data = 8'h00;
 2111 : data = 8'h00;
 2112 : data = 8'h00;
 2113 : data = 8'h00;
 2114 : data = 8'h00;
 2115 : data = 8'h00;
 2116 : data = 8'h00;
 2117 : data = 8'h00;
 2118 : data = 8'h00;
 2119 : data = 8'h00;
 2120 : data = 8'h00;
 2121 : data = 8'h00;
 2122 : data = 8'h00;
 2123 : data = 8'h00;
 2124 : data = 8'h00;
 2125 : data = 8'h00;
 2126 : data = 8'h00;
 2127 : data = 8'h00;
 2128 : data = 8'h00;
 2129 : data = 8'h00;
 2130 : data = 8'h00;
 2131 : data = 8'h00;
 2132 : data = 8'h00;
 2133 : data = 8'h00;
 2134 : data = 8'h00;
 2135 : data = 8'h00;
 2136 : data = 8'h00;
 2137 : data = 8'h00;
 2138 : data = 8'h00;
 2139 : data = 8'h00;
 2140 : data = 8'h00;
 2141 : data = 8'h00;
 2142 : data = 8'h00;
 2143 : data = 8'h00;
 2144 : data = 8'h00;
 2145 : data = 8'h00;
 2146 : data = 8'h00;
 2147 : data = 8'h00;
 2148 : data = 8'h00;
 2149 : data = 8'h00;
 2150 : data = 8'h00;
 2151 : data = 8'h00;
 2152 : data = 8'h00;
 2153 : data = 8'h00;
 2154 : data = 8'h00;
 2155 : data = 8'h00;
 2156 : data = 8'h00;
 2157 : data = 8'h00;
 2158 : data = 8'h00;
 2159 : data = 8'h00;
 2160 : data = 8'h00;
 2161 : data = 8'h00;
 2162 : data = 8'h00;
 2163 : data = 8'h00;
 2164 : data = 8'h00;
 2165 : data = 8'h00;
 2166 : data = 8'h00;
 2167 : data = 8'h00;
 2168 : data = 8'h00;
 2169 : data = 8'h00;
 2170 : data = 8'h00;
 2171 : data = 8'h00;
 2172 : data = 8'h00;
 2173 : data = 8'h00;
 2174 : data = 8'h00;
 2175 : data = 8'h00;
 2176 : data = 8'h00;
 2177 : data = 8'h00;
 2178 : data = 8'h00;
 2179 : data = 8'h00;
 2180 : data = 8'h00;
 2181 : data = 8'h00;
 2182 : data = 8'h00;
 2183 : data = 8'h00;
 2184 : data = 8'h00;
 2185 : data = 8'h00;
 2186 : data = 8'h00;
 2187 : data = 8'h00;
 2188 : data = 8'h00;
 2189 : data = 8'h00;
 2190 : data = 8'h00;
 2191 : data = 8'h00;
 2192 : data = 8'h00;
 2193 : data = 8'h00;
 2194 : data = 8'h00;
 2195 : data = 8'h00;
 2196 : data = 8'h00;
 2197 : data = 8'h00;
 2198 : data = 8'h00;
 2199 : data = 8'h00;
 2200 : data = 8'h00;
 2201 : data = 8'h00;
 2202 : data = 8'h00;
 2203 : data = 8'h00;
 2204 : data = 8'h00;
 2205 : data = 8'h00;
 2206 : data = 8'h00;
 2207 : data = 8'h00;
 2208 : data = 8'h00;
 2209 : data = 8'h00;
 2210 : data = 8'h00;
 2211 : data = 8'h00;
 2212 : data = 8'h00;
 2213 : data = 8'h00;
 2214 : data = 8'h00;
 2215 : data = 8'h00;
 2216 : data = 8'h00;
 2217 : data = 8'h00;
 2218 : data = 8'h00;
 2219 : data = 8'h00;
 2220 : data = 8'h00;
 2221 : data = 8'h00;
 2222 : data = 8'h00;
 2223 : data = 8'h00;
 2224 : data = 8'h00;
 2225 : data = 8'h00;
 2226 : data = 8'h00;
 2227 : data = 8'h00;
 2228 : data = 8'h00;
 2229 : data = 8'h00;
 2230 : data = 8'h00;
 2231 : data = 8'h00;
 2232 : data = 8'h00;
 2233 : data = 8'h00;
 2234 : data = 8'h00;
 2235 : data = 8'h00;
 2236 : data = 8'h00;
 2237 : data = 8'h00;
 2238 : data = 8'h00;
 2239 : data = 8'h00;
 2240 : data = 8'h00;
 2241 : data = 8'h00;
 2242 : data = 8'h00;
 2243 : data = 8'h00;
 2244 : data = 8'h00;
 2245 : data = 8'h00;
 2246 : data = 8'h00;
 2247 : data = 8'h00;
 2248 : data = 8'h00;
 2249 : data = 8'h00;
 2250 : data = 8'h00;
 2251 : data = 8'h00;
 2252 : data = 8'h00;
 2253 : data = 8'h00;
 2254 : data = 8'h00;
 2255 : data = 8'h00;
 2256 : data = 8'h00;
 2257 : data = 8'h00;
 2258 : data = 8'h00;
 2259 : data = 8'h00;
 2260 : data = 8'h00;
 2261 : data = 8'h00;
 2262 : data = 8'h00;
 2263 : data = 8'h00;
 2264 : data = 8'h00;
 2265 : data = 8'h00;
 2266 : data = 8'h00;
 2267 : data = 8'h00;
 2268 : data = 8'h00;
 2269 : data = 8'h00;
 2270 : data = 8'h00;
 2271 : data = 8'h00;
 2272 : data = 8'h00;
 2273 : data = 8'h00;
 2274 : data = 8'h00;
 2275 : data = 8'h00;
 2276 : data = 8'h00;
 2277 : data = 8'h00;
 2278 : data = 8'h00;
 2279 : data = 8'h00;
 2280 : data = 8'h00;
 2281 : data = 8'h00;
 2282 : data = 8'h00;
 2283 : data = 8'h00;
 2284 : data = 8'h00;
 2285 : data = 8'h00;
 2286 : data = 8'h00;
 2287 : data = 8'h00;
 2288 : data = 8'h00;
 2289 : data = 8'h00;
 2290 : data = 8'h00;
 2291 : data = 8'h00;
 2292 : data = 8'h00;
 2293 : data = 8'h00;
 2294 : data = 8'h00;
 2295 : data = 8'h00;
 2296 : data = 8'h00;
 2297 : data = 8'h00;
 2298 : data = 8'h00;
 2299 : data = 8'h00;
 2300 : data = 8'h00;
 2301 : data = 8'h00;
 2302 : data = 8'h00;
 2303 : data = 8'h00;
 2304 : data = 8'h00;
 2305 : data = 8'h00;
 2306 : data = 8'h00;
 2307 : data = 8'h00;
 2308 : data = 8'h00;
 2309 : data = 8'h00;
 2310 : data = 8'h00;
 2311 : data = 8'h00;
 2312 : data = 8'h00;
 2313 : data = 8'h00;
 2314 : data = 8'h00;
 2315 : data = 8'h00;
 2316 : data = 8'h00;
 2317 : data = 8'h00;
 2318 : data = 8'h00;
 2319 : data = 8'h00;
 2320 : data = 8'h00;
 2321 : data = 8'h00;
 2322 : data = 8'h00;
 2323 : data = 8'h00;
 2324 : data = 8'h00;
 2325 : data = 8'h00;
 2326 : data = 8'h00;
 2327 : data = 8'h00;
 2328 : data = 8'h00;
 2329 : data = 8'h00;
 2330 : data = 8'h00;
 2331 : data = 8'h00;
 2332 : data = 8'h00;
 2333 : data = 8'h00;
 2334 : data = 8'h00;
 2335 : data = 8'h00;
 2336 : data = 8'h00;
 2337 : data = 8'h00;
 2338 : data = 8'h00;
 2339 : data = 8'h00;
 2340 : data = 8'h00;
 2341 : data = 8'h00;
 2342 : data = 8'h00;
 2343 : data = 8'h00;
 2344 : data = 8'h00;
 2345 : data = 8'h00;
 2346 : data = 8'h00;
 2347 : data = 8'h00;
 2348 : data = 8'h00;
 2349 : data = 8'h00;
 2350 : data = 8'h00;
 2351 : data = 8'h00;
 2352 : data = 8'h00;
 2353 : data = 8'h00;
 2354 : data = 8'h00;
 2355 : data = 8'h00;
 2356 : data = 8'h00;
 2357 : data = 8'h00;
 2358 : data = 8'h00;
 2359 : data = 8'h00;
 2360 : data = 8'h00;
 2361 : data = 8'h00;
 2362 : data = 8'h00;
 2363 : data = 8'h00;
 2364 : data = 8'h00;
 2365 : data = 8'h00;
 2366 : data = 8'h00;
 2367 : data = 8'h00;
 2368 : data = 8'h00;
 2369 : data = 8'h00;
 2370 : data = 8'h00;
 2371 : data = 8'h00;
 2372 : data = 8'h00;
 2373 : data = 8'h00;
 2374 : data = 8'h00;
 2375 : data = 8'h00;
 2376 : data = 8'h00;
 2377 : data = 8'h00;
 2378 : data = 8'h00;
 2379 : data = 8'h00;
 2380 : data = 8'h00;
 2381 : data = 8'h00;
 2382 : data = 8'h00;
 2383 : data = 8'h00;
 2384 : data = 8'h00;
 2385 : data = 8'h00;
 2386 : data = 8'h00;
 2387 : data = 8'h00;
 2388 : data = 8'h00;
 2389 : data = 8'h00;
 2390 : data = 8'h00;
 2391 : data = 8'h00;
 2392 : data = 8'h00;
 2393 : data = 8'h00;
 2394 : data = 8'h00;
 2395 : data = 8'h00;
 2396 : data = 8'h00;
 2397 : data = 8'h00;
 2398 : data = 8'h00;
 2399 : data = 8'h00;
 2400 : data = 8'h00;
 2401 : data = 8'h00;
 2402 : data = 8'h00;
 2403 : data = 8'h00;
 2404 : data = 8'h00;
 2405 : data = 8'h00;
 2406 : data = 8'h00;
 2407 : data = 8'h00;
 2408 : data = 8'h00;
 2409 : data = 8'h00;
 2410 : data = 8'h00;
 2411 : data = 8'h00;
 2412 : data = 8'h00;
 2413 : data = 8'h00;
 2414 : data = 8'h00;
 2415 : data = 8'h00;
 2416 : data = 8'h00;
 2417 : data = 8'h00;
 2418 : data = 8'h00;
 2419 : data = 8'h00;
 2420 : data = 8'h00;
 2421 : data = 8'h00;
 2422 : data = 8'h00;
 2423 : data = 8'h00;
 2424 : data = 8'h00;
 2425 : data = 8'h00;
 2426 : data = 8'h00;
 2427 : data = 8'h00;
 2428 : data = 8'h00;
 2429 : data = 8'h00;
 2430 : data = 8'h00;
 2431 : data = 8'h00;
 2432 : data = 8'h00;
 2433 : data = 8'h00;
 2434 : data = 8'h00;
 2435 : data = 8'h00;
 2436 : data = 8'h00;
 2437 : data = 8'h00;
 2438 : data = 8'h00;
 2439 : data = 8'h00;
 2440 : data = 8'h00;
 2441 : data = 8'h00;
 2442 : data = 8'h00;
 2443 : data = 8'h00;
 2444 : data = 8'h00;
 2445 : data = 8'h00;
 2446 : data = 8'h00;
 2447 : data = 8'h00;
 2448 : data = 8'h00;
 2449 : data = 8'h00;
 2450 : data = 8'h00;
 2451 : data = 8'h00;
 2452 : data = 8'h00;
 2453 : data = 8'h00;
 2454 : data = 8'h00;
 2455 : data = 8'h00;
 2456 : data = 8'h00;
 2457 : data = 8'h00;
 2458 : data = 8'h00;
 2459 : data = 8'h00;
 2460 : data = 8'h00;
 2461 : data = 8'h00;
 2462 : data = 8'h00;
 2463 : data = 8'h00;
 2464 : data = 8'h00;
 2465 : data = 8'h00;
 2466 : data = 8'h00;
 2467 : data = 8'h00;
 2468 : data = 8'h00;
 2469 : data = 8'h00;
 2470 : data = 8'h00;
 2471 : data = 8'h00;
 2472 : data = 8'h00;
 2473 : data = 8'h00;
 2474 : data = 8'h00;
 2475 : data = 8'h00;
 2476 : data = 8'h00;
 2477 : data = 8'h00;
 2478 : data = 8'h00;
 2479 : data = 8'h00;
 2480 : data = 8'h00;
 2481 : data = 8'h00;
 2482 : data = 8'h00;
 2483 : data = 8'h00;
 2484 : data = 8'h00;
 2485 : data = 8'h00;
 2486 : data = 8'h00;
 2487 : data = 8'h00;
 2488 : data = 8'h00;
 2489 : data = 8'h00;
 2490 : data = 8'h00;
 2491 : data = 8'h00;
 2492 : data = 8'h00;
 2493 : data = 8'h00;
 2494 : data = 8'h00;
 2495 : data = 8'h00;
 2496 : data = 8'h00;
 2497 : data = 8'h00;
 2498 : data = 8'h00;
 2499 : data = 8'h00;
 2500 : data = 8'h00;
 2501 : data = 8'h00;
 2502 : data = 8'h00;
 2503 : data = 8'h00;
 2504 : data = 8'h00;
 2505 : data = 8'h00;
 2506 : data = 8'h00;
 2507 : data = 8'h00;
 2508 : data = 8'h00;
 2509 : data = 8'h00;
 2510 : data = 8'h00;
 2511 : data = 8'h00;
 2512 : data = 8'h00;
 2513 : data = 8'h00;
 2514 : data = 8'h00;
 2515 : data = 8'h00;
 2516 : data = 8'h00;
 2517 : data = 8'h00;
 2518 : data = 8'h00;
 2519 : data = 8'h00;
 2520 : data = 8'h00;
 2521 : data = 8'h00;
 2522 : data = 8'h00;
 2523 : data = 8'h00;
 2524 : data = 8'h00;
 2525 : data = 8'h00;
 2526 : data = 8'h00;
 2527 : data = 8'h00;
 2528 : data = 8'h00;
 2529 : data = 8'h00;
 2530 : data = 8'h00;
 2531 : data = 8'h00;
 2532 : data = 8'h00;
 2533 : data = 8'h00;
 2534 : data = 8'h00;
 2535 : data = 8'h00;
 2536 : data = 8'h00;
 2537 : data = 8'h00;
 2538 : data = 8'h00;
 2539 : data = 8'h00;
 2540 : data = 8'h00;
 2541 : data = 8'h00;
 2542 : data = 8'h00;
 2543 : data = 8'h00;
 2544 : data = 8'h00;
 2545 : data = 8'h00;
 2546 : data = 8'h00;
 2547 : data = 8'h00;
 2548 : data = 8'h00;
 2549 : data = 8'h00;
 2550 : data = 8'h00;
 2551 : data = 8'h00;
 2552 : data = 8'h00;
 2553 : data = 8'h00;
 2554 : data = 8'h00;
 2555 : data = 8'h00;
 2556 : data = 8'h00;
 2557 : data = 8'h00;
 2558 : data = 8'h00;
 2559 : data = 8'h00;
 2560 : data = 8'h00;
 2561 : data = 8'h00;
 2562 : data = 8'h00;
 2563 : data = 8'h00;
 2564 : data = 8'h00;
 2565 : data = 8'h00;
 2566 : data = 8'h00;
 2567 : data = 8'h00;
 2568 : data = 8'h00;
 2569 : data = 8'h00;
 2570 : data = 8'h00;
 2571 : data = 8'h00;
 2572 : data = 8'h00;
 2573 : data = 8'h00;
 2574 : data = 8'h00;
 2575 : data = 8'h00;
 2576 : data = 8'h00;
 2577 : data = 8'h00;
 2578 : data = 8'h00;
 2579 : data = 8'h00;
 2580 : data = 8'h00;
 2581 : data = 8'h00;
 2582 : data = 8'h00;
 2583 : data = 8'h00;
 2584 : data = 8'h00;
 2585 : data = 8'h00;
 2586 : data = 8'h00;
 2587 : data = 8'h00;
 2588 : data = 8'h00;
 2589 : data = 8'h00;
 2590 : data = 8'h00;
 2591 : data = 8'h00;
 2592 : data = 8'h00;
 2593 : data = 8'h00;
 2594 : data = 8'h00;
 2595 : data = 8'h00;
 2596 : data = 8'h00;
 2597 : data = 8'h00;
 2598 : data = 8'h00;
 2599 : data = 8'h00;
 2600 : data = 8'h00;
 2601 : data = 8'h00;
 2602 : data = 8'h00;
 2603 : data = 8'h00;
 2604 : data = 8'h00;
 2605 : data = 8'h00;
 2606 : data = 8'h00;
 2607 : data = 8'h00;
 2608 : data = 8'h00;
 2609 : data = 8'h00;
 2610 : data = 8'h00;
 2611 : data = 8'h00;
 2612 : data = 8'h00;
 2613 : data = 8'h00;
 2614 : data = 8'h00;
 2615 : data = 8'h00;
 2616 : data = 8'h00;
 2617 : data = 8'h00;
 2618 : data = 8'h00;
 2619 : data = 8'h00;
 2620 : data = 8'h00;
 2621 : data = 8'h00;
 2622 : data = 8'h00;
 2623 : data = 8'h00;
 2624 : data = 8'h00;
 2625 : data = 8'h00;
 2626 : data = 8'h00;
 2627 : data = 8'h00;
 2628 : data = 8'h00;
 2629 : data = 8'h00;
 2630 : data = 8'h00;
 2631 : data = 8'h00;
 2632 : data = 8'h00;
 2633 : data = 8'h00;
 2634 : data = 8'h00;
 2635 : data = 8'h00;
 2636 : data = 8'h00;
 2637 : data = 8'h00;
 2638 : data = 8'h00;
 2639 : data = 8'h00;
 2640 : data = 8'h00;
 2641 : data = 8'h00;
 2642 : data = 8'h00;
 2643 : data = 8'h00;
 2644 : data = 8'h00;
 2645 : data = 8'h00;
 2646 : data = 8'h00;
 2647 : data = 8'h00;
 2648 : data = 8'h00;
 2649 : data = 8'h00;
 2650 : data = 8'h00;
 2651 : data = 8'h00;
 2652 : data = 8'h00;
 2653 : data = 8'h00;
 2654 : data = 8'h00;
 2655 : data = 8'h00;
 2656 : data = 8'h00;
 2657 : data = 8'h00;
 2658 : data = 8'h00;
 2659 : data = 8'h00;
 2660 : data = 8'h00;
 2661 : data = 8'h00;
 2662 : data = 8'h00;
 2663 : data = 8'h00;
 2664 : data = 8'h00;
 2665 : data = 8'h00;
 2666 : data = 8'h00;
 2667 : data = 8'h00;
 2668 : data = 8'h00;
 2669 : data = 8'h00;
 2670 : data = 8'h00;
 2671 : data = 8'h00;
 2672 : data = 8'h00;
 2673 : data = 8'h00;
 2674 : data = 8'h00;
 2675 : data = 8'h00;
 2676 : data = 8'h00;
 2677 : data = 8'h00;
 2678 : data = 8'h00;
 2679 : data = 8'h00;
 2680 : data = 8'h00;
 2681 : data = 8'h00;
 2682 : data = 8'h00;
 2683 : data = 8'h00;
 2684 : data = 8'h00;
 2685 : data = 8'h00;
 2686 : data = 8'h00;
 2687 : data = 8'h00;
 2688 : data = 8'h00;
 2689 : data = 8'h00;
 2690 : data = 8'h00;
 2691 : data = 8'h00;
 2692 : data = 8'h00;
 2693 : data = 8'h00;
 2694 : data = 8'h00;
 2695 : data = 8'h00;
 2696 : data = 8'h00;
 2697 : data = 8'h00;
 2698 : data = 8'h00;
 2699 : data = 8'h00;
 2700 : data = 8'h00;
 2701 : data = 8'h00;
 2702 : data = 8'h00;
 2703 : data = 8'h00;
 2704 : data = 8'h00;
 2705 : data = 8'h00;
 2706 : data = 8'h00;
 2707 : data = 8'h00;
 2708 : data = 8'h00;
 2709 : data = 8'h00;
 2710 : data = 8'h00;
 2711 : data = 8'h00;
 2712 : data = 8'h00;
 2713 : data = 8'h00;
 2714 : data = 8'h00;
 2715 : data = 8'h00;
 2716 : data = 8'h00;
 2717 : data = 8'h00;
 2718 : data = 8'h00;
 2719 : data = 8'h00;
 2720 : data = 8'h00;
 2721 : data = 8'h00;
 2722 : data = 8'h00;
 2723 : data = 8'h00;
 2724 : data = 8'h00;
 2725 : data = 8'h00;
 2726 : data = 8'h00;
 2727 : data = 8'h00;
 2728 : data = 8'h00;
 2729 : data = 8'h00;
 2730 : data = 8'h00;
 2731 : data = 8'h00;
 2732 : data = 8'h00;
 2733 : data = 8'h00;
 2734 : data = 8'h00;
 2735 : data = 8'h00;
 2736 : data = 8'h00;
 2737 : data = 8'h00;
 2738 : data = 8'h00;
 2739 : data = 8'h00;
 2740 : data = 8'h00;
 2741 : data = 8'h00;
 2742 : data = 8'h00;
 2743 : data = 8'h00;
 2744 : data = 8'h00;
 2745 : data = 8'h00;
 2746 : data = 8'h00;
 2747 : data = 8'h00;
 2748 : data = 8'h00;
 2749 : data = 8'h00;
 2750 : data = 8'h00;
 2751 : data = 8'h00;
 2752 : data = 8'h00;
 2753 : data = 8'h00;
 2754 : data = 8'h00;
 2755 : data = 8'h00;
 2756 : data = 8'h00;
 2757 : data = 8'h00;
 2758 : data = 8'h00;
 2759 : data = 8'h00;
 2760 : data = 8'h00;
 2761 : data = 8'h00;
 2762 : data = 8'h00;
 2763 : data = 8'h00;
 2764 : data = 8'h00;
 2765 : data = 8'h00;
 2766 : data = 8'h00;
 2767 : data = 8'h00;
 2768 : data = 8'h00;
 2769 : data = 8'h00;
 2770 : data = 8'h00;
 2771 : data = 8'h00;
 2772 : data = 8'h00;
 2773 : data = 8'h00;
 2774 : data = 8'h00;
 2775 : data = 8'h00;
 2776 : data = 8'h00;
 2777 : data = 8'h00;
 2778 : data = 8'h00;
 2779 : data = 8'h00;
 2780 : data = 8'h00;
 2781 : data = 8'h00;
 2782 : data = 8'h00;
 2783 : data = 8'h00;
 2784 : data = 8'h00;
 2785 : data = 8'h00;
 2786 : data = 8'h00;
 2787 : data = 8'h00;
 2788 : data = 8'h00;
 2789 : data = 8'h00;
 2790 : data = 8'h00;
 2791 : data = 8'h00;
 2792 : data = 8'h00;
 2793 : data = 8'h00;
 2794 : data = 8'h00;
 2795 : data = 8'h00;
 2796 : data = 8'h00;
 2797 : data = 8'h00;
 2798 : data = 8'h00;
 2799 : data = 8'h00;
 2800 : data = 8'h00;
 2801 : data = 8'h00;
 2802 : data = 8'h00;
 2803 : data = 8'h00;
 2804 : data = 8'h00;
 2805 : data = 8'h00;
 2806 : data = 8'h00;
 2807 : data = 8'h00;
 2808 : data = 8'h00;
 2809 : data = 8'h00;
 2810 : data = 8'h00;
 2811 : data = 8'h00;
 2812 : data = 8'h00;
 2813 : data = 8'h00;
 2814 : data = 8'h00;
 2815 : data = 8'h00;
 2816 : data = 8'h00;
 2817 : data = 8'h00;
 2818 : data = 8'h00;
 2819 : data = 8'h00;
 2820 : data = 8'h00;
 2821 : data = 8'h00;
 2822 : data = 8'h00;
 2823 : data = 8'h00;
 2824 : data = 8'h00;
 2825 : data = 8'h00;
 2826 : data = 8'h00;
 2827 : data = 8'h00;
 2828 : data = 8'h00;
 2829 : data = 8'h00;
 2830 : data = 8'h00;
 2831 : data = 8'h00;
 2832 : data = 8'h00;
 2833 : data = 8'h00;
 2834 : data = 8'h00;
 2835 : data = 8'h00;
 2836 : data = 8'h00;
 2837 : data = 8'h00;
 2838 : data = 8'h00;
 2839 : data = 8'h00;
 2840 : data = 8'h00;
 2841 : data = 8'h00;
 2842 : data = 8'h00;
 2843 : data = 8'h00;
 2844 : data = 8'h00;
 2845 : data = 8'h00;
 2846 : data = 8'h00;
 2847 : data = 8'h00;
 2848 : data = 8'h00;
 2849 : data = 8'h00;
 2850 : data = 8'h00;
 2851 : data = 8'h00;
 2852 : data = 8'h00;
 2853 : data = 8'h00;
 2854 : data = 8'h00;
 2855 : data = 8'h00;
 2856 : data = 8'h00;
 2857 : data = 8'h00;
 2858 : data = 8'h00;
 2859 : data = 8'h00;
 2860 : data = 8'h00;
 2861 : data = 8'h00;
 2862 : data = 8'h00;
 2863 : data = 8'h00;
 2864 : data = 8'h00;
 2865 : data = 8'h00;
 2866 : data = 8'h00;
 2867 : data = 8'h00;
 2868 : data = 8'h00;
 2869 : data = 8'h00;
 2870 : data = 8'h00;
 2871 : data = 8'h00;
 2872 : data = 8'h00;
 2873 : data = 8'h00;
 2874 : data = 8'h00;
 2875 : data = 8'h00;
 2876 : data = 8'h00;
 2877 : data = 8'h00;
 2878 : data = 8'h00;
 2879 : data = 8'h00;
 2880 : data = 8'h00;
 2881 : data = 8'h00;
 2882 : data = 8'h00;
 2883 : data = 8'h00;
 2884 : data = 8'h00;
 2885 : data = 8'h00;
 2886 : data = 8'h00;
 2887 : data = 8'h00;
 2888 : data = 8'h00;
 2889 : data = 8'h00;
 2890 : data = 8'h00;
 2891 : data = 8'h00;
 2892 : data = 8'h00;
 2893 : data = 8'h00;
 2894 : data = 8'h00;
 2895 : data = 8'h00;
 2896 : data = 8'h00;
 2897 : data = 8'h00;
 2898 : data = 8'h00;
 2899 : data = 8'h00;
 2900 : data = 8'h00;
 2901 : data = 8'h00;
 2902 : data = 8'h00;
 2903 : data = 8'h00;
 2904 : data = 8'h00;
 2905 : data = 8'h00;
 2906 : data = 8'h00;
 2907 : data = 8'h00;
 2908 : data = 8'h00;
 2909 : data = 8'h00;
 2910 : data = 8'h00;
 2911 : data = 8'h00;
 2912 : data = 8'h00;
 2913 : data = 8'h00;
 2914 : data = 8'h00;
 2915 : data = 8'h00;
 2916 : data = 8'h00;
 2917 : data = 8'h00;
 2918 : data = 8'h00;
 2919 : data = 8'h00;
 2920 : data = 8'h00;
 2921 : data = 8'h00;
 2922 : data = 8'h00;
 2923 : data = 8'h00;
 2924 : data = 8'h00;
 2925 : data = 8'h00;
 2926 : data = 8'h00;
 2927 : data = 8'h00;
 2928 : data = 8'h00;
 2929 : data = 8'h00;
 2930 : data = 8'h00;
 2931 : data = 8'h00;
 2932 : data = 8'h00;
 2933 : data = 8'h00;
 2934 : data = 8'h00;
 2935 : data = 8'h00;
 2936 : data = 8'h00;
 2937 : data = 8'h00;
 2938 : data = 8'h00;
 2939 : data = 8'h00;
 2940 : data = 8'h00;
 2941 : data = 8'h00;
 2942 : data = 8'h00;
 2943 : data = 8'h00;
 2944 : data = 8'h00;
 2945 : data = 8'h00;
 2946 : data = 8'h00;
 2947 : data = 8'h00;
 2948 : data = 8'h00;
 2949 : data = 8'h00;
 2950 : data = 8'h00;
 2951 : data = 8'h00;
 2952 : data = 8'h00;
 2953 : data = 8'h00;
 2954 : data = 8'h00;
 2955 : data = 8'h00;
 2956 : data = 8'h00;
 2957 : data = 8'h00;
 2958 : data = 8'h00;
 2959 : data = 8'h00;
 2960 : data = 8'h00;
 2961 : data = 8'h00;
 2962 : data = 8'h00;
 2963 : data = 8'h00;
 2964 : data = 8'h00;
 2965 : data = 8'h00;
 2966 : data = 8'h00;
 2967 : data = 8'h00;
 2968 : data = 8'h00;
 2969 : data = 8'h00;
 2970 : data = 8'h00;
 2971 : data = 8'h00;
 2972 : data = 8'h00;
 2973 : data = 8'h00;
 2974 : data = 8'h00;
 2975 : data = 8'h00;
 2976 : data = 8'h00;
 2977 : data = 8'h00;
 2978 : data = 8'h00;
 2979 : data = 8'h00;
 2980 : data = 8'h00;
 2981 : data = 8'h00;
 2982 : data = 8'h00;
 2983 : data = 8'h00;
 2984 : data = 8'h00;
 2985 : data = 8'h00;
 2986 : data = 8'h00;
 2987 : data = 8'h00;
 2988 : data = 8'h00;
 2989 : data = 8'h00;
 2990 : data = 8'h00;
 2991 : data = 8'h00;
 2992 : data = 8'h00;
 2993 : data = 8'h00;
 2994 : data = 8'h00;
 2995 : data = 8'h00;
 2996 : data = 8'h00;
 2997 : data = 8'h00;
 2998 : data = 8'h00;
 2999 : data = 8'h00;
 3000 : data = 8'h00;
 3001 : data = 8'h00;
 3002 : data = 8'h00;
 3003 : data = 8'h00;
 3004 : data = 8'h00;
 3005 : data = 8'h00;
 3006 : data = 8'h00;
 3007 : data = 8'h00;
 3008 : data = 8'h00;
 3009 : data = 8'h00;
 3010 : data = 8'h00;
 3011 : data = 8'h00;
 3012 : data = 8'h00;
 3013 : data = 8'h00;
 3014 : data = 8'h00;
 3015 : data = 8'h00;
 3016 : data = 8'h00;
 3017 : data = 8'h00;
 3018 : data = 8'h00;
 3019 : data = 8'h00;
 3020 : data = 8'h00;
 3021 : data = 8'h00;
 3022 : data = 8'h00;
 3023 : data = 8'h00;
 3024 : data = 8'h00;
 3025 : data = 8'h00;
 3026 : data = 8'h00;
 3027 : data = 8'h00;
 3028 : data = 8'h00;
 3029 : data = 8'h00;
 3030 : data = 8'h00;
 3031 : data = 8'h00;
 3032 : data = 8'h00;
 3033 : data = 8'h00;
 3034 : data = 8'h00;
 3035 : data = 8'h00;
 3036 : data = 8'h00;
 3037 : data = 8'h00;
 3038 : data = 8'h00;
 3039 : data = 8'h00;
 3040 : data = 8'h00;
 3041 : data = 8'h00;
 3042 : data = 8'h00;
 3043 : data = 8'h00;
 3044 : data = 8'h00;
 3045 : data = 8'h00;
 3046 : data = 8'h00;
 3047 : data = 8'h00;
 3048 : data = 8'h00;
 3049 : data = 8'h00;
 3050 : data = 8'h00;
 3051 : data = 8'h00;
 3052 : data = 8'h00;
 3053 : data = 8'h00;
 3054 : data = 8'h00;
 3055 : data = 8'h00;
 3056 : data = 8'h00;
 3057 : data = 8'h00;
 3058 : data = 8'h00;
 3059 : data = 8'h00;
 3060 : data = 8'h00;
 3061 : data = 8'h00;
 3062 : data = 8'h00;
 3063 : data = 8'h00;
 3064 : data = 8'h00;
 3065 : data = 8'h00;
 3066 : data = 8'h00;
 3067 : data = 8'h00;
 3068 : data = 8'h00;
 3069 : data = 8'h00;
 3070 : data = 8'h00;
 3071 : data = 8'h00;
 3072 : data = 8'h00;
 3073 : data = 8'h00;
 3074 : data = 8'h00;
 3075 : data = 8'h00;
 3076 : data = 8'h00;
 3077 : data = 8'h00;
 3078 : data = 8'h00;
 3079 : data = 8'h00;
 3080 : data = 8'h00;
 3081 : data = 8'h00;
 3082 : data = 8'h00;
 3083 : data = 8'h00;
 3084 : data = 8'h00;
 3085 : data = 8'h00;
 3086 : data = 8'h00;
 3087 : data = 8'h00;
 3088 : data = 8'h00;
 3089 : data = 8'h00;
 3090 : data = 8'h00;
 3091 : data = 8'h00;
 3092 : data = 8'h00;
 3093 : data = 8'h00;
 3094 : data = 8'h00;
 3095 : data = 8'h00;
 3096 : data = 8'h00;
 3097 : data = 8'h00;
 3098 : data = 8'h00;
 3099 : data = 8'h00;
 3100 : data = 8'h00;
 3101 : data = 8'h00;
 3102 : data = 8'h00;
 3103 : data = 8'h00;
 3104 : data = 8'h00;
 3105 : data = 8'h00;
 3106 : data = 8'h00;
 3107 : data = 8'h00;
 3108 : data = 8'h00;
 3109 : data = 8'h00;
 3110 : data = 8'h00;
 3111 : data = 8'h00;
 3112 : data = 8'h00;
 3113 : data = 8'h00;
 3114 : data = 8'h00;
 3115 : data = 8'h00;
 3116 : data = 8'h00;
 3117 : data = 8'h00;
 3118 : data = 8'h00;
 3119 : data = 8'h00;
 3120 : data = 8'h00;
 3121 : data = 8'h00;
 3122 : data = 8'h00;
 3123 : data = 8'h00;
 3124 : data = 8'h00;
 3125 : data = 8'h00;
 3126 : data = 8'h00;
 3127 : data = 8'h00;
 3128 : data = 8'h00;
 3129 : data = 8'h00;
 3130 : data = 8'h00;
 3131 : data = 8'h00;
 3132 : data = 8'h00;
 3133 : data = 8'h00;
 3134 : data = 8'h00;
 3135 : data = 8'h00;
 3136 : data = 8'h00;
 3137 : data = 8'h00;
 3138 : data = 8'h00;
 3139 : data = 8'h00;
 3140 : data = 8'h00;
 3141 : data = 8'h00;
 3142 : data = 8'h00;
 3143 : data = 8'h00;
 3144 : data = 8'h00;
 3145 : data = 8'h00;
 3146 : data = 8'h00;
 3147 : data = 8'h00;
 3148 : data = 8'h00;
 3149 : data = 8'h00;
 3150 : data = 8'h00;
 3151 : data = 8'h00;
 3152 : data = 8'h00;
 3153 : data = 8'h00;
 3154 : data = 8'h00;
 3155 : data = 8'h00;
 3156 : data = 8'h00;
 3157 : data = 8'h00;
 3158 : data = 8'h00;
 3159 : data = 8'h00;
 3160 : data = 8'h00;
 3161 : data = 8'h00;
 3162 : data = 8'h00;
 3163 : data = 8'h00;
 3164 : data = 8'h00;
 3165 : data = 8'h00;
 3166 : data = 8'h00;
 3167 : data = 8'h00;
 3168 : data = 8'h00;
 3169 : data = 8'h00;
 3170 : data = 8'h00;
 3171 : data = 8'h00;
 3172 : data = 8'h00;
 3173 : data = 8'h00;
 3174 : data = 8'h00;
 3175 : data = 8'h00;
 3176 : data = 8'h00;
 3177 : data = 8'h00;
 3178 : data = 8'h00;
 3179 : data = 8'h00;
 3180 : data = 8'h00;
 3181 : data = 8'h00;
 3182 : data = 8'h00;
 3183 : data = 8'h00;
 3184 : data = 8'h00;
 3185 : data = 8'h00;
 3186 : data = 8'h00;
 3187 : data = 8'h00;
 3188 : data = 8'h00;
 3189 : data = 8'h00;
 3190 : data = 8'h00;
 3191 : data = 8'h00;
 3192 : data = 8'h00;
 3193 : data = 8'h00;
 3194 : data = 8'h00;
 3195 : data = 8'h00;
 3196 : data = 8'h00;
 3197 : data = 8'h00;
 3198 : data = 8'h00;
 3199 : data = 8'h00;
 3200 : data = 8'h00;
 3201 : data = 8'h00;
 3202 : data = 8'h00;
 3203 : data = 8'h00;
 3204 : data = 8'h00;
 3205 : data = 8'h00;
 3206 : data = 8'h00;
 3207 : data = 8'h00;
 3208 : data = 8'h00;
 3209 : data = 8'h00;
 3210 : data = 8'h00;
 3211 : data = 8'h00;
 3212 : data = 8'h00;
 3213 : data = 8'h00;
 3214 : data = 8'h00;
 3215 : data = 8'h00;
 3216 : data = 8'h00;
 3217 : data = 8'h00;
 3218 : data = 8'h00;
 3219 : data = 8'h00;
 3220 : data = 8'h00;
 3221 : data = 8'h00;
 3222 : data = 8'h00;
 3223 : data = 8'h00;
 3224 : data = 8'h00;
 3225 : data = 8'h00;
 3226 : data = 8'h00;
 3227 : data = 8'h00;
 3228 : data = 8'h00;
 3229 : data = 8'h00;
 3230 : data = 8'h00;
 3231 : data = 8'h00;
 3232 : data = 8'h00;
 3233 : data = 8'h00;
 3234 : data = 8'h00;
 3235 : data = 8'h00;
 3236 : data = 8'h00;
 3237 : data = 8'h00;
 3238 : data = 8'h00;
 3239 : data = 8'h00;
 3240 : data = 8'h00;
 3241 : data = 8'h00;
 3242 : data = 8'h00;
 3243 : data = 8'h00;
 3244 : data = 8'h00;
 3245 : data = 8'h00;
 3246 : data = 8'h00;
 3247 : data = 8'h00;
 3248 : data = 8'h00;
 3249 : data = 8'h00;
 3250 : data = 8'h00;
 3251 : data = 8'h00;
 3252 : data = 8'h00;
 3253 : data = 8'h00;
 3254 : data = 8'h00;
 3255 : data = 8'h00;
 3256 : data = 8'h00;
 3257 : data = 8'h00;
 3258 : data = 8'h00;
 3259 : data = 8'h00;
 3260 : data = 8'h00;
 3261 : data = 8'h00;
 3262 : data = 8'h00;
 3263 : data = 8'h00;
 3264 : data = 8'h00;
 3265 : data = 8'h00;
 3266 : data = 8'h00;
 3267 : data = 8'h00;
 3268 : data = 8'h00;
 3269 : data = 8'h00;
 3270 : data = 8'h00;
 3271 : data = 8'h00;
 3272 : data = 8'h00;
 3273 : data = 8'h00;
 3274 : data = 8'h00;
 3275 : data = 8'h00;
 3276 : data = 8'h00;
 3277 : data = 8'h00;
 3278 : data = 8'h00;
 3279 : data = 8'h00;
 3280 : data = 8'h00;
 3281 : data = 8'h00;
 3282 : data = 8'h00;
 3283 : data = 8'h00;
 3284 : data = 8'h00;
 3285 : data = 8'h00;
 3286 : data = 8'h00;
 3287 : data = 8'h00;
 3288 : data = 8'h00;
 3289 : data = 8'h00;
 3290 : data = 8'h00;
 3291 : data = 8'h00;
 3292 : data = 8'h00;
 3293 : data = 8'h00;
 3294 : data = 8'h00;
 3295 : data = 8'h00;
 3296 : data = 8'h00;
 3297 : data = 8'h00;
 3298 : data = 8'h00;
 3299 : data = 8'h00;
 3300 : data = 8'h00;
 3301 : data = 8'h00;
 3302 : data = 8'h00;
 3303 : data = 8'h00;
 3304 : data = 8'h00;
 3305 : data = 8'h00;
 3306 : data = 8'h00;
 3307 : data = 8'h00;
 3308 : data = 8'h00;
 3309 : data = 8'h00;
 3310 : data = 8'h00;
 3311 : data = 8'h00;
 3312 : data = 8'h00;
 3313 : data = 8'h00;
 3314 : data = 8'h00;
 3315 : data = 8'h00;
 3316 : data = 8'h00;
 3317 : data = 8'h00;
 3318 : data = 8'h00;
 3319 : data = 8'h00;
 3320 : data = 8'h00;
 3321 : data = 8'h00;
 3322 : data = 8'h00;
 3323 : data = 8'h00;
 3324 : data = 8'h00;
 3325 : data = 8'h00;
 3326 : data = 8'h00;
 3327 : data = 8'h00;
 3328 : data = 8'h00;
 3329 : data = 8'h00;
 3330 : data = 8'h00;
 3331 : data = 8'h00;
 3332 : data = 8'h00;
 3333 : data = 8'h00;
 3334 : data = 8'h00;
 3335 : data = 8'h00;
 3336 : data = 8'h00;
 3337 : data = 8'h00;
 3338 : data = 8'h00;
 3339 : data = 8'h00;
 3340 : data = 8'h00;
 3341 : data = 8'h00;
 3342 : data = 8'h00;
 3343 : data = 8'h00;
 3344 : data = 8'h00;
 3345 : data = 8'h00;
 3346 : data = 8'h00;
 3347 : data = 8'h00;
 3348 : data = 8'h00;
 3349 : data = 8'h00;
 3350 : data = 8'h00;
 3351 : data = 8'h00;
 3352 : data = 8'h00;
 3353 : data = 8'h00;
 3354 : data = 8'h00;
 3355 : data = 8'h00;
 3356 : data = 8'h00;
 3357 : data = 8'h00;
 3358 : data = 8'h00;
 3359 : data = 8'h00;
 3360 : data = 8'h00;
 3361 : data = 8'h00;
 3362 : data = 8'h00;
 3363 : data = 8'h00;
 3364 : data = 8'h00;
 3365 : data = 8'h00;
 3366 : data = 8'h00;
 3367 : data = 8'h00;
 3368 : data = 8'h00;
 3369 : data = 8'h00;
 3370 : data = 8'h00;
 3371 : data = 8'h00;
 3372 : data = 8'h00;
 3373 : data = 8'h00;
 3374 : data = 8'h00;
 3375 : data = 8'h00;
 3376 : data = 8'h00;
 3377 : data = 8'h00;
 3378 : data = 8'h00;
 3379 : data = 8'h00;
 3380 : data = 8'h00;
 3381 : data = 8'h00;
 3382 : data = 8'h00;
 3383 : data = 8'h00;
 3384 : data = 8'h00;
 3385 : data = 8'h00;
 3386 : data = 8'h00;
 3387 : data = 8'h00;
 3388 : data = 8'h00;
 3389 : data = 8'h00;
 3390 : data = 8'h00;
 3391 : data = 8'h00;
 3392 : data = 8'h00;
 3393 : data = 8'h00;
 3394 : data = 8'h00;
 3395 : data = 8'h00;
 3396 : data = 8'h00;
 3397 : data = 8'h00;
 3398 : data = 8'h00;
 3399 : data = 8'h00;
 3400 : data = 8'h00;
 3401 : data = 8'h00;
 3402 : data = 8'h00;
 3403 : data = 8'h00;
 3404 : data = 8'h00;
 3405 : data = 8'h00;
 3406 : data = 8'h00;
 3407 : data = 8'h00;
 3408 : data = 8'h00;
 3409 : data = 8'h00;
 3410 : data = 8'h00;
 3411 : data = 8'h00;
 3412 : data = 8'h00;
 3413 : data = 8'h00;
 3414 : data = 8'h00;
 3415 : data = 8'h00;
 3416 : data = 8'h00;
 3417 : data = 8'h00;
 3418 : data = 8'h00;
 3419 : data = 8'h00;
 3420 : data = 8'h00;
 3421 : data = 8'h00;
 3422 : data = 8'h00;
 3423 : data = 8'h00;
 3424 : data = 8'h00;
 3425 : data = 8'h00;
 3426 : data = 8'h00;
 3427 : data = 8'h00;
 3428 : data = 8'h00;
 3429 : data = 8'h00;
 3430 : data = 8'h00;
 3431 : data = 8'h00;
 3432 : data = 8'h00;
 3433 : data = 8'h00;
 3434 : data = 8'h00;
 3435 : data = 8'h00;
 3436 : data = 8'h00;
 3437 : data = 8'h00;
 3438 : data = 8'h00;
 3439 : data = 8'h00;
 3440 : data = 8'h00;
 3441 : data = 8'h00;
 3442 : data = 8'h00;
 3443 : data = 8'h00;
 3444 : data = 8'h00;
 3445 : data = 8'h00;
 3446 : data = 8'h00;
 3447 : data = 8'h00;
 3448 : data = 8'h00;
 3449 : data = 8'h00;
 3450 : data = 8'h00;
 3451 : data = 8'h00;
 3452 : data = 8'h00;
 3453 : data = 8'h00;
 3454 : data = 8'h00;
 3455 : data = 8'h00;
 3456 : data = 8'h00;
 3457 : data = 8'h00;
 3458 : data = 8'h00;
 3459 : data = 8'h00;
 3460 : data = 8'h00;
 3461 : data = 8'h00;
 3462 : data = 8'h00;
 3463 : data = 8'h00;
 3464 : data = 8'h00;
 3465 : data = 8'h00;
 3466 : data = 8'h00;
 3467 : data = 8'h00;
 3468 : data = 8'h00;
 3469 : data = 8'h00;
 3470 : data = 8'h00;
 3471 : data = 8'h00;
 3472 : data = 8'h00;
 3473 : data = 8'h00;
 3474 : data = 8'h00;
 3475 : data = 8'h00;
 3476 : data = 8'h00;
 3477 : data = 8'h00;
 3478 : data = 8'h00;
 3479 : data = 8'h00;
 3480 : data = 8'h00;
 3481 : data = 8'h00;
 3482 : data = 8'h00;
 3483 : data = 8'h00;
 3484 : data = 8'h00;
 3485 : data = 8'h00;
 3486 : data = 8'h00;
 3487 : data = 8'h00;
 3488 : data = 8'h00;
 3489 : data = 8'h00;
 3490 : data = 8'h00;
 3491 : data = 8'h00;
 3492 : data = 8'h00;
 3493 : data = 8'h00;
 3494 : data = 8'h00;
 3495 : data = 8'h00;
 3496 : data = 8'h00;
 3497 : data = 8'h00;
 3498 : data = 8'h00;
 3499 : data = 8'h00;
 3500 : data = 8'h00;
 3501 : data = 8'h00;
 3502 : data = 8'h00;
 3503 : data = 8'h00;
 3504 : data = 8'h00;
 3505 : data = 8'h00;
 3506 : data = 8'h00;
 3507 : data = 8'h00;
 3508 : data = 8'h00;
 3509 : data = 8'h00;
 3510 : data = 8'h00;
 3511 : data = 8'h00;
 3512 : data = 8'h00;
 3513 : data = 8'h00;
 3514 : data = 8'h00;
 3515 : data = 8'h00;
 3516 : data = 8'h00;
 3517 : data = 8'h00;
 3518 : data = 8'h00;
 3519 : data = 8'h00;
 3520 : data = 8'h00;
 3521 : data = 8'h00;
 3522 : data = 8'h00;
 3523 : data = 8'h00;
 3524 : data = 8'h00;
 3525 : data = 8'h00;
 3526 : data = 8'h00;
 3527 : data = 8'h00;
 3528 : data = 8'h00;
 3529 : data = 8'h00;
 3530 : data = 8'h00;
 3531 : data = 8'h00;
 3532 : data = 8'h00;
 3533 : data = 8'h00;
 3534 : data = 8'h00;
 3535 : data = 8'h00;
 3536 : data = 8'h00;
 3537 : data = 8'h00;
 3538 : data = 8'h00;
 3539 : data = 8'h00;
 3540 : data = 8'h00;
 3541 : data = 8'h00;
 3542 : data = 8'h00;
 3543 : data = 8'h00;
 3544 : data = 8'h00;
 3545 : data = 8'h00;
 3546 : data = 8'h00;
 3547 : data = 8'h00;
 3548 : data = 8'h00;
 3549 : data = 8'h00;
 3550 : data = 8'h00;
 3551 : data = 8'h00;
 3552 : data = 8'h00;
 3553 : data = 8'h00;
 3554 : data = 8'h00;
 3555 : data = 8'h00;
 3556 : data = 8'h00;
 3557 : data = 8'h00;
 3558 : data = 8'h00;
 3559 : data = 8'h00;
 3560 : data = 8'h00;
 3561 : data = 8'h00;
 3562 : data = 8'h00;
 3563 : data = 8'h00;
 3564 : data = 8'h00;
 3565 : data = 8'h00;
 3566 : data = 8'h00;
 3567 : data = 8'h00;
 3568 : data = 8'h00;
 3569 : data = 8'h00;
 3570 : data = 8'h00;
 3571 : data = 8'h00;
 3572 : data = 8'h00;
 3573 : data = 8'h00;
 3574 : data = 8'h00;
 3575 : data = 8'h00;
 3576 : data = 8'h00;
 3577 : data = 8'h00;
 3578 : data = 8'h00;
 3579 : data = 8'h00;
 3580 : data = 8'h00;
 3581 : data = 8'h00;
 3582 : data = 8'h00;
 3583 : data = 8'h00;
 3584 : data = 8'h00;
 3585 : data = 8'h00;
 3586 : data = 8'h00;
 3587 : data = 8'h00;
 3588 : data = 8'h00;
 3589 : data = 8'h00;
 3590 : data = 8'h00;
 3591 : data = 8'h00;
 3592 : data = 8'h00;
 3593 : data = 8'h00;
 3594 : data = 8'h00;
 3595 : data = 8'h00;
 3596 : data = 8'h00;
 3597 : data = 8'h00;
 3598 : data = 8'h00;
 3599 : data = 8'h00;
 3600 : data = 8'h00;
 3601 : data = 8'h00;
 3602 : data = 8'h00;
 3603 : data = 8'h00;
 3604 : data = 8'h00;
 3605 : data = 8'h00;
 3606 : data = 8'h00;
 3607 : data = 8'h00;
 3608 : data = 8'h00;
 3609 : data = 8'h00;
 3610 : data = 8'h00;
 3611 : data = 8'h00;
 3612 : data = 8'h00;
 3613 : data = 8'h00;
 3614 : data = 8'h00;
 3615 : data = 8'h00;
 3616 : data = 8'h00;
 3617 : data = 8'h00;
 3618 : data = 8'h00;
 3619 : data = 8'h00;
 3620 : data = 8'h00;
 3621 : data = 8'h00;
 3622 : data = 8'h00;
 3623 : data = 8'h00;
 3624 : data = 8'h00;
 3625 : data = 8'h00;
 3626 : data = 8'h00;
 3627 : data = 8'h00;
 3628 : data = 8'h00;
 3629 : data = 8'h00;
 3630 : data = 8'h00;
 3631 : data = 8'h00;
 3632 : data = 8'h00;
 3633 : data = 8'h00;
 3634 : data = 8'h00;
 3635 : data = 8'h00;
 3636 : data = 8'h00;
 3637 : data = 8'h00;
 3638 : data = 8'h00;
 3639 : data = 8'h00;
 3640 : data = 8'h00;
 3641 : data = 8'h00;
 3642 : data = 8'h00;
 3643 : data = 8'h00;
 3644 : data = 8'h00;
 3645 : data = 8'h00;
 3646 : data = 8'h00;
 3647 : data = 8'h00;
 3648 : data = 8'h00;
 3649 : data = 8'h00;
 3650 : data = 8'h00;
 3651 : data = 8'h00;
 3652 : data = 8'h00;
 3653 : data = 8'h00;
 3654 : data = 8'h00;
 3655 : data = 8'h00;
 3656 : data = 8'h00;
 3657 : data = 8'h00;
 3658 : data = 8'h00;
 3659 : data = 8'h00;
 3660 : data = 8'h00;
 3661 : data = 8'h00;
 3662 : data = 8'h00;
 3663 : data = 8'h00;
 3664 : data = 8'h00;
 3665 : data = 8'h00;
 3666 : data = 8'h00;
 3667 : data = 8'h00;
 3668 : data = 8'h00;
 3669 : data = 8'h00;
 3670 : data = 8'h00;
 3671 : data = 8'h00;
 3672 : data = 8'h00;
 3673 : data = 8'h00;
 3674 : data = 8'h00;
 3675 : data = 8'h00;
 3676 : data = 8'h00;
 3677 : data = 8'h00;
 3678 : data = 8'h00;
 3679 : data = 8'h00;
 3680 : data = 8'h00;
 3681 : data = 8'h00;
 3682 : data = 8'h00;
 3683 : data = 8'h00;
 3684 : data = 8'h00;
 3685 : data = 8'h00;
 3686 : data = 8'h00;
 3687 : data = 8'h00;
 3688 : data = 8'h00;
 3689 : data = 8'h00;
 3690 : data = 8'h00;
 3691 : data = 8'h00;
 3692 : data = 8'h00;
 3693 : data = 8'h00;
 3694 : data = 8'h00;
 3695 : data = 8'h00;
 3696 : data = 8'h00;
 3697 : data = 8'h00;
 3698 : data = 8'h00;
 3699 : data = 8'h00;
 3700 : data = 8'h00;
 3701 : data = 8'h00;
 3702 : data = 8'h00;
 3703 : data = 8'h00;
 3704 : data = 8'h00;
 3705 : data = 8'h00;
 3706 : data = 8'h00;
 3707 : data = 8'h00;
 3708 : data = 8'h00;
 3709 : data = 8'h00;
 3710 : data = 8'h00;
 3711 : data = 8'h00;
 3712 : data = 8'h00;
 3713 : data = 8'h00;
 3714 : data = 8'h00;
 3715 : data = 8'h00;
 3716 : data = 8'h00;
 3717 : data = 8'h00;
 3718 : data = 8'h00;
 3719 : data = 8'h00;
 3720 : data = 8'h00;
 3721 : data = 8'h00;
 3722 : data = 8'h00;
 3723 : data = 8'h00;
 3724 : data = 8'h00;
 3725 : data = 8'h00;
 3726 : data = 8'h00;
 3727 : data = 8'h00;
 3728 : data = 8'h00;
 3729 : data = 8'h00;
 3730 : data = 8'h00;
 3731 : data = 8'h00;
 3732 : data = 8'h00;
 3733 : data = 8'h00;
 3734 : data = 8'h00;
 3735 : data = 8'h00;
 3736 : data = 8'h00;
 3737 : data = 8'h00;
 3738 : data = 8'h00;
 3739 : data = 8'h00;
 3740 : data = 8'h00;
 3741 : data = 8'h00;
 3742 : data = 8'h00;
 3743 : data = 8'h00;
 3744 : data = 8'h00;
 3745 : data = 8'h00;
 3746 : data = 8'h00;
 3747 : data = 8'h00;
 3748 : data = 8'h00;
 3749 : data = 8'h00;
 3750 : data = 8'h00;
 3751 : data = 8'h00;
 3752 : data = 8'h00;
 3753 : data = 8'h00;
 3754 : data = 8'h00;
 3755 : data = 8'h00;
 3756 : data = 8'h00;
 3757 : data = 8'h00;
 3758 : data = 8'h00;
 3759 : data = 8'h00;
 3760 : data = 8'h00;
 3761 : data = 8'h00;
 3762 : data = 8'h00;
 3763 : data = 8'h00;
 3764 : data = 8'h00;
 3765 : data = 8'h00;
 3766 : data = 8'h00;
 3767 : data = 8'h00;
 3768 : data = 8'h00;
 3769 : data = 8'h00;
 3770 : data = 8'h00;
 3771 : data = 8'h00;
 3772 : data = 8'h00;
 3773 : data = 8'h00;
 3774 : data = 8'h00;
 3775 : data = 8'h00;
 3776 : data = 8'h00;
 3777 : data = 8'h00;
 3778 : data = 8'h00;
 3779 : data = 8'h00;
 3780 : data = 8'h00;
 3781 : data = 8'h00;
 3782 : data = 8'h00;
 3783 : data = 8'h00;
 3784 : data = 8'h00;
 3785 : data = 8'h00;
 3786 : data = 8'h00;
 3787 : data = 8'h00;
 3788 : data = 8'h00;
 3789 : data = 8'h00;
 3790 : data = 8'h00;
 3791 : data = 8'h00;
 3792 : data = 8'h00;
 3793 : data = 8'h00;
 3794 : data = 8'h00;
 3795 : data = 8'h00;
 3796 : data = 8'h00;
 3797 : data = 8'h00;
 3798 : data = 8'h00;
 3799 : data = 8'h00;
 3800 : data = 8'h00;
 3801 : data = 8'h00;
 3802 : data = 8'h00;
 3803 : data = 8'h00;
 3804 : data = 8'h00;
 3805 : data = 8'h00;
 3806 : data = 8'h00;
 3807 : data = 8'h00;
 3808 : data = 8'h00;
 3809 : data = 8'h00;
 3810 : data = 8'h00;
 3811 : data = 8'h00;
 3812 : data = 8'h00;
 3813 : data = 8'h00;
 3814 : data = 8'h00;
 3815 : data = 8'h00;
 3816 : data = 8'h00;
 3817 : data = 8'h00;
 3818 : data = 8'h00;
 3819 : data = 8'h00;
 3820 : data = 8'h00;
 3821 : data = 8'h00;
 3822 : data = 8'h00;
 3823 : data = 8'h00;
 3824 : data = 8'h00;
 3825 : data = 8'h00;
 3826 : data = 8'h00;
 3827 : data = 8'h00;
 3828 : data = 8'h00;
 3829 : data = 8'h00;
 3830 : data = 8'h00;
 3831 : data = 8'h00;
 3832 : data = 8'h00;
 3833 : data = 8'h00;
 3834 : data = 8'h00;
 3835 : data = 8'h00;
 3836 : data = 8'h00;
 3837 : data = 8'h00;
 3838 : data = 8'h00;
 3839 : data = 8'h00;
 3840 : data = 8'h00;
 3841 : data = 8'h00;
 3842 : data = 8'h00;
 3843 : data = 8'h00;
 3844 : data = 8'h00;
 3845 : data = 8'h00;
 3846 : data = 8'h00;
 3847 : data = 8'h00;
 3848 : data = 8'h00;
 3849 : data = 8'h00;
 3850 : data = 8'h00;
 3851 : data = 8'h00;
 3852 : data = 8'h00;
 3853 : data = 8'h00;
 3854 : data = 8'h00;
 3855 : data = 8'h00;
 3856 : data = 8'h00;
 3857 : data = 8'h00;
 3858 : data = 8'h00;
 3859 : data = 8'h00;
 3860 : data = 8'h00;
 3861 : data = 8'h00;
 3862 : data = 8'h00;
 3863 : data = 8'h00;
 3864 : data = 8'h00;
 3865 : data = 8'h00;
 3866 : data = 8'h00;
 3867 : data = 8'h00;
 3868 : data = 8'h00;
 3869 : data = 8'h00;
 3870 : data = 8'h00;
 3871 : data = 8'h00;
 3872 : data = 8'h00;
 3873 : data = 8'h00;
 3874 : data = 8'h00;
 3875 : data = 8'h00;
 3876 : data = 8'h00;
 3877 : data = 8'h00;
 3878 : data = 8'h00;
 3879 : data = 8'h00;
 3880 : data = 8'h00;
 3881 : data = 8'h00;
 3882 : data = 8'h00;
 3883 : data = 8'h00;
 3884 : data = 8'h00;
 3885 : data = 8'h00;
 3886 : data = 8'h00;
 3887 : data = 8'h00;
 3888 : data = 8'h00;
 3889 : data = 8'h00;
 3890 : data = 8'h00;
 3891 : data = 8'h00;
 3892 : data = 8'h00;
 3893 : data = 8'h00;
 3894 : data = 8'h00;
 3895 : data = 8'h00;
 3896 : data = 8'h00;
 3897 : data = 8'h00;
 3898 : data = 8'h00;
 3899 : data = 8'h00;
 3900 : data = 8'h00;
 3901 : data = 8'h00;
 3902 : data = 8'h00;
 3903 : data = 8'h00;
 3904 : data = 8'h00;
 3905 : data = 8'h00;
 3906 : data = 8'h00;
 3907 : data = 8'h00;
 3908 : data = 8'h00;
 3909 : data = 8'h00;
 3910 : data = 8'h00;
 3911 : data = 8'h00;
 3912 : data = 8'h00;
 3913 : data = 8'h00;
 3914 : data = 8'h00;
 3915 : data = 8'h00;
 3916 : data = 8'h00;
 3917 : data = 8'h00;
 3918 : data = 8'h00;
 3919 : data = 8'h00;
 3920 : data = 8'h00;
 3921 : data = 8'h00;
 3922 : data = 8'h00;
 3923 : data = 8'h00;
 3924 : data = 8'h00;
 3925 : data = 8'h00;
 3926 : data = 8'h00;
 3927 : data = 8'h00;
 3928 : data = 8'h00;
 3929 : data = 8'h00;
 3930 : data = 8'h00;
 3931 : data = 8'h00;
 3932 : data = 8'h00;
 3933 : data = 8'h00;
 3934 : data = 8'h00;
 3935 : data = 8'h00;
 3936 : data = 8'h00;
 3937 : data = 8'h00;
 3938 : data = 8'h00;
 3939 : data = 8'h00;
 3940 : data = 8'h00;
 3941 : data = 8'h00;
 3942 : data = 8'h00;
 3943 : data = 8'h00;
 3944 : data = 8'h00;
 3945 : data = 8'h00;
 3946 : data = 8'h00;
 3947 : data = 8'h00;
 3948 : data = 8'h00;
 3949 : data = 8'h00;
 3950 : data = 8'h00;
 3951 : data = 8'h00;
 3952 : data = 8'h00;
 3953 : data = 8'h00;
 3954 : data = 8'h00;
 3955 : data = 8'h00;
 3956 : data = 8'h00;
 3957 : data = 8'h00;
 3958 : data = 8'h00;
 3959 : data = 8'h00;
 3960 : data = 8'h00;
 3961 : data = 8'h00;
 3962 : data = 8'h00;
 3963 : data = 8'h00;
 3964 : data = 8'h00;
 3965 : data = 8'h00;
 3966 : data = 8'h00;
 3967 : data = 8'h00;
 3968 : data = 8'h00;
 3969 : data = 8'h00;
 3970 : data = 8'h00;
 3971 : data = 8'h00;
 3972 : data = 8'h00;
 3973 : data = 8'h00;
 3974 : data = 8'h00;
 3975 : data = 8'h00;
 3976 : data = 8'h00;
 3977 : data = 8'h00;
 3978 : data = 8'h00;
 3979 : data = 8'h00;
 3980 : data = 8'h00;
 3981 : data = 8'h00;
 3982 : data = 8'h00;
 3983 : data = 8'h00;
 3984 : data = 8'h00;
 3985 : data = 8'h00;
 3986 : data = 8'h00;
 3987 : data = 8'h00;
 3988 : data = 8'h00;
 3989 : data = 8'h00;
 3990 : data = 8'h00;
 3991 : data = 8'h00;
 3992 : data = 8'h00;
 3993 : data = 8'h00;
 3994 : data = 8'h00;
 3995 : data = 8'h00;
 3996 : data = 8'h00;
 3997 : data = 8'h00;
 3998 : data = 8'h00;
 3999 : data = 8'h00;
 4000 : data = 8'h00;
 4001 : data = 8'h00;
 4002 : data = 8'h00;
 4003 : data = 8'h00;
 4004 : data = 8'h00;
 4005 : data = 8'h00;
 4006 : data = 8'h00;
 4007 : data = 8'h00;
 4008 : data = 8'h00;
 4009 : data = 8'h00;
 4010 : data = 8'h00;
 4011 : data = 8'h00;
 4012 : data = 8'h00;
 4013 : data = 8'h00;
 4014 : data = 8'h00;
 4015 : data = 8'h00;
 4016 : data = 8'h00;
 4017 : data = 8'h00;
 4018 : data = 8'h00;
 4019 : data = 8'h00;
 4020 : data = 8'h00;
 4021 : data = 8'h00;
 4022 : data = 8'h00;
 4023 : data = 8'h00;
 4024 : data = 8'h00;
 4025 : data = 8'h00;
 4026 : data = 8'h00;
 4027 : data = 8'h00;
 4028 : data = 8'h00;
 4029 : data = 8'h00;
 4030 : data = 8'h00;
 4031 : data = 8'h00;
 4032 : data = 8'h00;
 4033 : data = 8'h00;
 4034 : data = 8'h00;
 4035 : data = 8'h00;
 4036 : data = 8'h00;
 4037 : data = 8'h00;
 4038 : data = 8'h00;
 4039 : data = 8'h00;
 4040 : data = 8'h00;
 4041 : data = 8'h00;
 4042 : data = 8'h00;
 4043 : data = 8'h00;
 4044 : data = 8'h00;
 4045 : data = 8'h00;
 4046 : data = 8'h00;
 4047 : data = 8'h00;
 4048 : data = 8'h00;
 4049 : data = 8'h00;
 4050 : data = 8'h00;
 4051 : data = 8'h00;
 4052 : data = 8'h00;
 4053 : data = 8'h00;
 4054 : data = 8'h00;
 4055 : data = 8'h00;
 4056 : data = 8'h00;
 4057 : data = 8'h00;
 4058 : data = 8'h00;
 4059 : data = 8'h00;
 4060 : data = 8'h00;
 4061 : data = 8'h00;
 4062 : data = 8'h00;
 4063 : data = 8'h00;
 4064 : data = 8'h00;
 4065 : data = 8'h00;
 4066 : data = 8'h00;
 4067 : data = 8'h00;
 4068 : data = 8'h00;
 4069 : data = 8'h00;
 4070 : data = 8'h00;
 4071 : data = 8'h00;
 4072 : data = 8'h00;
 4073 : data = 8'h00;
 4074 : data = 8'h00;
 4075 : data = 8'h00;
 4076 : data = 8'h00;
 4077 : data = 8'h00;
 4078 : data = 8'h00;
 4079 : data = 8'h00;
 4080 : data = 8'h00;
 4081 : data = 8'h00;
 4082 : data = 8'h00;
 4083 : data = 8'h00;
 4084 : data = 8'h00;
 4085 : data = 8'h00;
 4086 : data = 8'h00;
 4087 : data = 8'h00;
 4088 : data = 8'h00;
 4089 : data = 8'h00;
 4090 : data = 8'h00;
 4091 : data = 8'h00;
 4092 : data = 8'h00;
 4093 : data = 8'h00;
 4094 : data = 8'h00;
 4095 : data = 8'h00;
 4096 : data = 8'h00;
 4097 : data = 8'h00;
 4098 : data = 8'h00;
 4099 : data = 8'h00;
 4100 : data = 8'h00;
 4101 : data = 8'h00;
 4102 : data = 8'h00;
 4103 : data = 8'h00;
 4104 : data = 8'h00;
 4105 : data = 8'h00;
 4106 : data = 8'h00;
 4107 : data = 8'h00;
 4108 : data = 8'h00;
 4109 : data = 8'h00;
 4110 : data = 8'h00;
 4111 : data = 8'h00;
 4112 : data = 8'h00;
 4113 : data = 8'h00;
 4114 : data = 8'h00;
 4115 : data = 8'h00;
 4116 : data = 8'h00;
 4117 : data = 8'h00;
 4118 : data = 8'h00;
 4119 : data = 8'h00;
 4120 : data = 8'h00;
 4121 : data = 8'h00;
 4122 : data = 8'h00;
 4123 : data = 8'h00;
 4124 : data = 8'h00;
 4125 : data = 8'h00;
 4126 : data = 8'h00;
 4127 : data = 8'h00;
 4128 : data = 8'h00;
 4129 : data = 8'h00;
 4130 : data = 8'h00;
 4131 : data = 8'h00;
 4132 : data = 8'h00;
 4133 : data = 8'h00;
 4134 : data = 8'h00;
 4135 : data = 8'h00;
 4136 : data = 8'h00;
 4137 : data = 8'h00;
 4138 : data = 8'h00;
 4139 : data = 8'h00;
 4140 : data = 8'h00;
 4141 : data = 8'h00;
 4142 : data = 8'h00;
 4143 : data = 8'h00;
 4144 : data = 8'h00;
 4145 : data = 8'h00;
 4146 : data = 8'h00;
 4147 : data = 8'h00;
 4148 : data = 8'h00;
 4149 : data = 8'h00;
 4150 : data = 8'h00;
 4151 : data = 8'h00;
 4152 : data = 8'h00;
 4153 : data = 8'h00;
 4154 : data = 8'h00;
 4155 : data = 8'h00;
 4156 : data = 8'h00;
 4157 : data = 8'h00;
 4158 : data = 8'h00;
 4159 : data = 8'h00;
 4160 : data = 8'h00;
 4161 : data = 8'h00;
 4162 : data = 8'h00;
 4163 : data = 8'h00;
 4164 : data = 8'h00;
 4165 : data = 8'h00;
 4166 : data = 8'h00;
 4167 : data = 8'h00;
 4168 : data = 8'h00;
 4169 : data = 8'h00;
 4170 : data = 8'h00;
 4171 : data = 8'h00;
 4172 : data = 8'h00;
 4173 : data = 8'h00;
 4174 : data = 8'h00;
 4175 : data = 8'h00;
 4176 : data = 8'h00;
 4177 : data = 8'h00;
 4178 : data = 8'h00;
 4179 : data = 8'h00;
 4180 : data = 8'h00;
 4181 : data = 8'h00;
 4182 : data = 8'h00;
 4183 : data = 8'h00;
 4184 : data = 8'h00;
 4185 : data = 8'h00;
 4186 : data = 8'h00;
 4187 : data = 8'h00;
 4188 : data = 8'h00;
 4189 : data = 8'h00;
 4190 : data = 8'h00;
 4191 : data = 8'h00;
 4192 : data = 8'h00;
 4193 : data = 8'h00;
 4194 : data = 8'h00;
 4195 : data = 8'h00;
 4196 : data = 8'h00;
 4197 : data = 8'h00;
 4198 : data = 8'h00;
 4199 : data = 8'h00;
 4200 : data = 8'h00;
 4201 : data = 8'h00;
 4202 : data = 8'h00;
 4203 : data = 8'h00;
 4204 : data = 8'h00;
 4205 : data = 8'h00;
 4206 : data = 8'h00;
 4207 : data = 8'h00;
 4208 : data = 8'h00;
 4209 : data = 8'h00;
 4210 : data = 8'h00;
 4211 : data = 8'h00;
 4212 : data = 8'h00;
 4213 : data = 8'h00;
 4214 : data = 8'h00;
 4215 : data = 8'h00;
 4216 : data = 8'h00;
 4217 : data = 8'h00;
 4218 : data = 8'h00;
 4219 : data = 8'h00;
 4220 : data = 8'h00;
 4221 : data = 8'h00;
 4222 : data = 8'h00;
 4223 : data = 8'h00;
 4224 : data = 8'h00;
 4225 : data = 8'h00;
 4226 : data = 8'h00;
 4227 : data = 8'h00;
 4228 : data = 8'h00;
 4229 : data = 8'h00;
 4230 : data = 8'h00;
 4231 : data = 8'h00;
 4232 : data = 8'h00;
 4233 : data = 8'h00;
 4234 : data = 8'h00;
 4235 : data = 8'h00;
 4236 : data = 8'h00;
 4237 : data = 8'h00;
 4238 : data = 8'h00;
 4239 : data = 8'h00;
 4240 : data = 8'h00;
 4241 : data = 8'h00;
 4242 : data = 8'h00;
 4243 : data = 8'h00;
 4244 : data = 8'h00;
 4245 : data = 8'h00;
 4246 : data = 8'h00;
 4247 : data = 8'h00;
 4248 : data = 8'h00;
 4249 : data = 8'h00;
 4250 : data = 8'h00;
 4251 : data = 8'h00;
 4252 : data = 8'h00;
 4253 : data = 8'h00;
 4254 : data = 8'h00;
 4255 : data = 8'h00;
 4256 : data = 8'h00;
 4257 : data = 8'h00;
 4258 : data = 8'h00;
 4259 : data = 8'h00;
 4260 : data = 8'h00;
 4261 : data = 8'h00;
 4262 : data = 8'h00;
 4263 : data = 8'h00;
 4264 : data = 8'h00;
 4265 : data = 8'h00;
 4266 : data = 8'h00;
 4267 : data = 8'h00;
 4268 : data = 8'h00;
 4269 : data = 8'h00;
 4270 : data = 8'h00;
 4271 : data = 8'h00;
 4272 : data = 8'h00;
 4273 : data = 8'h00;
 4274 : data = 8'h00;
 4275 : data = 8'h00;
 4276 : data = 8'h00;
 4277 : data = 8'h00;
 4278 : data = 8'h00;
 4279 : data = 8'h00;
 4280 : data = 8'h00;
 4281 : data = 8'h00;
 4282 : data = 8'h00;
 4283 : data = 8'h00;
 4284 : data = 8'h00;
 4285 : data = 8'h00;
 4286 : data = 8'h00;
 4287 : data = 8'h00;
 4288 : data = 8'h00;
 4289 : data = 8'h00;
 4290 : data = 8'h00;
 4291 : data = 8'h00;
 4292 : data = 8'h00;
 4293 : data = 8'h00;
 4294 : data = 8'h00;
 4295 : data = 8'h00;
 4296 : data = 8'h00;
 4297 : data = 8'h00;
 4298 : data = 8'h00;
 4299 : data = 8'h00;
 4300 : data = 8'h00;
 4301 : data = 8'h00;
 4302 : data = 8'h00;
 4303 : data = 8'h00;
 4304 : data = 8'h00;
 4305 : data = 8'h00;
 4306 : data = 8'h00;
 4307 : data = 8'h00;
 4308 : data = 8'h00;
 4309 : data = 8'h00;
 4310 : data = 8'h00;
 4311 : data = 8'h00;
 4312 : data = 8'h00;
 4313 : data = 8'h00;
 4314 : data = 8'h00;
 4315 : data = 8'h00;
 4316 : data = 8'h00;
 4317 : data = 8'h00;
 4318 : data = 8'h00;
 4319 : data = 8'h00;
 4320 : data = 8'h00;
 4321 : data = 8'h00;
 4322 : data = 8'h00;
 4323 : data = 8'h00;
 4324 : data = 8'h00;
 4325 : data = 8'h00;
 4326 : data = 8'h00;
 4327 : data = 8'h00;
 4328 : data = 8'h00;
 4329 : data = 8'h00;
 4330 : data = 8'h00;
 4331 : data = 8'h00;
 4332 : data = 8'h00;
 4333 : data = 8'h00;
 4334 : data = 8'h00;
 4335 : data = 8'h00;
 4336 : data = 8'h00;
 4337 : data = 8'h00;
 4338 : data = 8'h00;
 4339 : data = 8'h00;
 4340 : data = 8'h00;
 4341 : data = 8'h00;
 4342 : data = 8'h00;
 4343 : data = 8'h00;
 4344 : data = 8'h00;
 4345 : data = 8'h00;
 4346 : data = 8'h00;
 4347 : data = 8'h00;
 4348 : data = 8'h00;
 4349 : data = 8'h00;
 4350 : data = 8'h00;
 4351 : data = 8'h00;
 4352 : data = 8'h00;
 4353 : data = 8'h00;
 4354 : data = 8'h00;
 4355 : data = 8'h00;
 4356 : data = 8'h00;
 4357 : data = 8'h00;
 4358 : data = 8'h00;
 4359 : data = 8'h00;
 4360 : data = 8'h00;
 4361 : data = 8'h00;
 4362 : data = 8'h00;
 4363 : data = 8'h00;
 4364 : data = 8'h00;
 4365 : data = 8'h00;
 4366 : data = 8'h00;
 4367 : data = 8'h00;
 4368 : data = 8'h00;
 4369 : data = 8'h00;
 4370 : data = 8'h00;
 4371 : data = 8'h00;
 4372 : data = 8'h00;
 4373 : data = 8'h00;
 4374 : data = 8'h00;
 4375 : data = 8'h00;
 4376 : data = 8'h00;
 4377 : data = 8'h00;
 4378 : data = 8'h00;
 4379 : data = 8'h00;
 4380 : data = 8'h00;
 4381 : data = 8'h00;
 4382 : data = 8'h00;
 4383 : data = 8'h00;
 4384 : data = 8'h00;
 4385 : data = 8'h00;
 4386 : data = 8'h00;
 4387 : data = 8'h00;
 4388 : data = 8'h00;
 4389 : data = 8'h00;
 4390 : data = 8'h00;
 4391 : data = 8'h00;
 4392 : data = 8'h00;
 4393 : data = 8'h00;
 4394 : data = 8'h00;
 4395 : data = 8'h00;
 4396 : data = 8'h00;
 4397 : data = 8'h00;
 4398 : data = 8'h00;
 4399 : data = 8'h00;
 4400 : data = 8'h00;
 4401 : data = 8'h00;
 4402 : data = 8'h00;
 4403 : data = 8'h00;
 4404 : data = 8'h00;
 4405 : data = 8'h00;
 4406 : data = 8'h00;
 4407 : data = 8'h00;
 4408 : data = 8'h00;
 4409 : data = 8'h00;
 4410 : data = 8'h00;
 4411 : data = 8'h00;
 4412 : data = 8'h00;
 4413 : data = 8'h00;
 4414 : data = 8'h00;
 4415 : data = 8'h00;
 4416 : data = 8'h00;
 4417 : data = 8'h00;
 4418 : data = 8'h00;
 4419 : data = 8'h00;
 4420 : data = 8'h00;
 4421 : data = 8'h00;
 4422 : data = 8'h00;
 4423 : data = 8'h00;
 4424 : data = 8'h00;
 4425 : data = 8'h00;
 4426 : data = 8'h00;
 4427 : data = 8'h00;
 4428 : data = 8'h00;
 4429 : data = 8'h00;
 4430 : data = 8'h00;
 4431 : data = 8'h00;
 4432 : data = 8'h00;
 4433 : data = 8'h00;
 4434 : data = 8'h00;
 4435 : data = 8'h00;
 4436 : data = 8'h00;
 4437 : data = 8'h00;
 4438 : data = 8'h00;
 4439 : data = 8'h00;
 4440 : data = 8'h00;
 4441 : data = 8'h00;
 4442 : data = 8'h00;
 4443 : data = 8'h00;
 4444 : data = 8'h00;
 4445 : data = 8'h00;
 4446 : data = 8'h00;
 4447 : data = 8'h00;
 4448 : data = 8'h00;
 4449 : data = 8'h00;
 4450 : data = 8'h00;
 4451 : data = 8'h00;
 4452 : data = 8'h00;
 4453 : data = 8'h00;
 4454 : data = 8'h00;
 4455 : data = 8'h00;
 4456 : data = 8'h00;
 4457 : data = 8'h00;
 4458 : data = 8'h00;
 4459 : data = 8'h00;
 4460 : data = 8'h00;
 4461 : data = 8'h00;
 4462 : data = 8'h00;
 4463 : data = 8'h00;
 4464 : data = 8'h00;
 4465 : data = 8'h00;
 4466 : data = 8'h00;
 4467 : data = 8'h00;
 4468 : data = 8'h00;
 4469 : data = 8'h00;
 4470 : data = 8'h00;
 4471 : data = 8'h00;
 4472 : data = 8'h00;
 4473 : data = 8'h00;
 4474 : data = 8'h00;
 4475 : data = 8'h00;
 4476 : data = 8'h00;
 4477 : data = 8'h00;
 4478 : data = 8'h00;
 4479 : data = 8'h00;
 4480 : data = 8'h00;
 4481 : data = 8'h00;
 4482 : data = 8'h00;
 4483 : data = 8'h00;
 4484 : data = 8'h00;
 4485 : data = 8'h00;
 4486 : data = 8'h00;
 4487 : data = 8'h00;
 4488 : data = 8'h00;
 4489 : data = 8'h00;
 4490 : data = 8'h00;
 4491 : data = 8'h00;
 4492 : data = 8'h00;
 4493 : data = 8'h00;
 4494 : data = 8'h00;
 4495 : data = 8'h00;
 4496 : data = 8'h00;
 4497 : data = 8'h00;
 4498 : data = 8'h00;
 4499 : data = 8'h00;
 4500 : data = 8'h00;
 4501 : data = 8'h00;
 4502 : data = 8'h00;
 4503 : data = 8'h00;
 4504 : data = 8'h00;
 4505 : data = 8'h00;
 4506 : data = 8'h00;
 4507 : data = 8'h00;
 4508 : data = 8'h00;
 4509 : data = 8'h00;
 4510 : data = 8'h00;
 4511 : data = 8'h00;
 4512 : data = 8'h00;
 4513 : data = 8'h00;
 4514 : data = 8'h00;
 4515 : data = 8'h00;
 4516 : data = 8'h00;
 4517 : data = 8'h00;
 4518 : data = 8'h00;
 4519 : data = 8'h00;
 4520 : data = 8'h00;
 4521 : data = 8'h00;
 4522 : data = 8'h00;
 4523 : data = 8'h00;
 4524 : data = 8'h00;
 4525 : data = 8'h00;
 4526 : data = 8'h00;
 4527 : data = 8'h00;
 4528 : data = 8'h00;
 4529 : data = 8'h00;
 4530 : data = 8'h00;
 4531 : data = 8'h00;
 4532 : data = 8'h00;
 4533 : data = 8'h00;
 4534 : data = 8'h00;
 4535 : data = 8'h00;
 4536 : data = 8'h00;
 4537 : data = 8'h00;
 4538 : data = 8'h00;
 4539 : data = 8'h00;
 4540 : data = 8'h00;
 4541 : data = 8'h00;
 4542 : data = 8'h00;
 4543 : data = 8'h00;
 4544 : data = 8'h00;
 4545 : data = 8'h00;
 4546 : data = 8'h00;
 4547 : data = 8'h00;
 4548 : data = 8'h00;
 4549 : data = 8'h00;
 4550 : data = 8'h00;
 4551 : data = 8'h00;
 4552 : data = 8'h00;
 4553 : data = 8'h00;
 4554 : data = 8'h00;
 4555 : data = 8'h00;
 4556 : data = 8'h00;
 4557 : data = 8'h00;
 4558 : data = 8'h00;
 4559 : data = 8'h00;
 4560 : data = 8'h00;
 4561 : data = 8'h00;
 4562 : data = 8'h00;
 4563 : data = 8'h00;
 4564 : data = 8'h00;
 4565 : data = 8'h00;
 4566 : data = 8'h00;
 4567 : data = 8'h00;
 4568 : data = 8'h00;
 4569 : data = 8'h00;
 4570 : data = 8'h00;
 4571 : data = 8'h00;
 4572 : data = 8'h00;
 4573 : data = 8'h00;
 4574 : data = 8'h00;
 4575 : data = 8'h00;
 4576 : data = 8'h00;
 4577 : data = 8'h00;
 4578 : data = 8'h00;
 4579 : data = 8'h00;
 4580 : data = 8'h00;
 4581 : data = 8'h00;
 4582 : data = 8'h00;
 4583 : data = 8'h00;
 4584 : data = 8'h00;
 4585 : data = 8'h00;
 4586 : data = 8'h00;
 4587 : data = 8'h00;
 4588 : data = 8'h00;
 4589 : data = 8'h00;
 4590 : data = 8'h00;
 4591 : data = 8'h00;
 4592 : data = 8'h00;
 4593 : data = 8'h00;
 4594 : data = 8'h00;
 4595 : data = 8'h00;
 4596 : data = 8'h00;
 4597 : data = 8'h00;
 4598 : data = 8'h00;
 4599 : data = 8'h00;
 4600 : data = 8'h00;
 4601 : data = 8'h00;
 4602 : data = 8'h00;
 4603 : data = 8'h00;
 4604 : data = 8'h00;
 4605 : data = 8'h00;
 4606 : data = 8'h00;
 4607 : data = 8'h00;
 4608 : data = 8'h00;
 4609 : data = 8'h00;
 4610 : data = 8'h00;
 4611 : data = 8'h00;
 4612 : data = 8'h00;
 4613 : data = 8'h00;
 4614 : data = 8'h00;
 4615 : data = 8'h00;
 4616 : data = 8'h00;
 4617 : data = 8'h00;
 4618 : data = 8'h00;
 4619 : data = 8'h00;
 4620 : data = 8'h00;
 4621 : data = 8'h00;
 4622 : data = 8'h00;
 4623 : data = 8'h00;
 4624 : data = 8'h00;
 4625 : data = 8'h00;
 4626 : data = 8'h00;
 4627 : data = 8'h00;
 4628 : data = 8'h00;
 4629 : data = 8'h00;
 4630 : data = 8'h00;
 4631 : data = 8'h00;
 4632 : data = 8'h00;
 4633 : data = 8'h00;
 4634 : data = 8'h00;
 4635 : data = 8'h00;
 4636 : data = 8'h00;
 4637 : data = 8'h00;
 4638 : data = 8'h00;
 4639 : data = 8'h00;
 4640 : data = 8'h00;
 4641 : data = 8'h00;
 4642 : data = 8'h00;
 4643 : data = 8'h00;
 4644 : data = 8'h00;
 4645 : data = 8'h00;
 4646 : data = 8'h00;
 4647 : data = 8'h00;
 4648 : data = 8'h00;
 4649 : data = 8'h00;
 4650 : data = 8'h00;
 4651 : data = 8'h00;
 4652 : data = 8'h00;
 4653 : data = 8'h00;
 4654 : data = 8'h00;
 4655 : data = 8'h00;
 4656 : data = 8'h00;
 4657 : data = 8'h00;
 4658 : data = 8'h00;
 4659 : data = 8'h00;
 4660 : data = 8'h00;
 4661 : data = 8'h00;
 4662 : data = 8'h00;
 4663 : data = 8'h00;
 4664 : data = 8'h00;
 4665 : data = 8'h00;
 4666 : data = 8'h00;
 4667 : data = 8'h00;
 4668 : data = 8'h00;
 4669 : data = 8'h00;
 4670 : data = 8'h00;
 4671 : data = 8'h00;
 4672 : data = 8'h00;
 4673 : data = 8'h00;
 4674 : data = 8'h00;
 4675 : data = 8'h00;
 4676 : data = 8'h00;
 4677 : data = 8'h00;
 4678 : data = 8'h00;
 4679 : data = 8'h00;
 4680 : data = 8'h00;
 4681 : data = 8'h00;
 4682 : data = 8'h00;
 4683 : data = 8'h00;
 4684 : data = 8'h00;
 4685 : data = 8'h00;
 4686 : data = 8'h00;
 4687 : data = 8'h00;
 4688 : data = 8'h00;
 4689 : data = 8'h00;
 4690 : data = 8'h00;
 4691 : data = 8'h00;
 4692 : data = 8'h00;
 4693 : data = 8'h00;
 4694 : data = 8'h00;
 4695 : data = 8'h00;
 4696 : data = 8'h00;
 4697 : data = 8'h00;
 4698 : data = 8'h00;
 4699 : data = 8'h00;
 4700 : data = 8'h00;
 4701 : data = 8'h00;
 4702 : data = 8'h00;
 4703 : data = 8'h00;
 4704 : data = 8'h00;
 4705 : data = 8'h00;
 4706 : data = 8'h00;
 4707 : data = 8'h00;
 4708 : data = 8'h00;
 4709 : data = 8'h00;
 4710 : data = 8'h00;
 4711 : data = 8'h00;
 4712 : data = 8'h00;
 4713 : data = 8'h00;
 4714 : data = 8'h00;
 4715 : data = 8'h00;
 4716 : data = 8'h00;
 4717 : data = 8'h00;
 4718 : data = 8'h00;
 4719 : data = 8'h00;
 4720 : data = 8'h00;
 4721 : data = 8'h00;
 4722 : data = 8'h00;
 4723 : data = 8'h00;
 4724 : data = 8'h00;
 4725 : data = 8'h00;
 4726 : data = 8'h00;
 4727 : data = 8'h00;
 4728 : data = 8'h00;
 4729 : data = 8'h00;
 4730 : data = 8'h00;
 4731 : data = 8'h00;
 4732 : data = 8'h00;
 4733 : data = 8'h00;
 4734 : data = 8'h00;
 4735 : data = 8'h00;
 4736 : data = 8'h00;
 4737 : data = 8'h00;
 4738 : data = 8'h00;
 4739 : data = 8'h00;
 4740 : data = 8'h00;
 4741 : data = 8'h00;
 4742 : data = 8'h00;
 4743 : data = 8'h00;
 4744 : data = 8'h00;
 4745 : data = 8'h00;
 4746 : data = 8'h00;
 4747 : data = 8'h00;
 4748 : data = 8'h00;
 4749 : data = 8'h00;
 4750 : data = 8'h00;
 4751 : data = 8'h00;
 4752 : data = 8'h00;
 4753 : data = 8'h00;
 4754 : data = 8'h00;
 4755 : data = 8'h00;
 4756 : data = 8'h00;
 4757 : data = 8'h00;
 4758 : data = 8'h00;
 4759 : data = 8'h00;
 4760 : data = 8'h00;
 4761 : data = 8'h00;
 4762 : data = 8'h00;
 4763 : data = 8'h00;
 4764 : data = 8'h00;
 4765 : data = 8'h00;
 4766 : data = 8'h00;
 4767 : data = 8'h00;
 4768 : data = 8'h00;
 4769 : data = 8'h00;
 4770 : data = 8'h00;
 4771 : data = 8'h00;
 4772 : data = 8'h00;
 4773 : data = 8'h00;
 4774 : data = 8'h00;
 4775 : data = 8'h00;
 4776 : data = 8'h00;
 4777 : data = 8'h00;
 4778 : data = 8'h00;
 4779 : data = 8'h00;
 4780 : data = 8'h00;
 4781 : data = 8'h00;
 4782 : data = 8'h00;
 4783 : data = 8'h00;
 4784 : data = 8'h00;
 4785 : data = 8'h00;
 4786 : data = 8'h00;
 4787 : data = 8'h00;
 4788 : data = 8'h00;
 4789 : data = 8'h00;
 4790 : data = 8'h00;
 4791 : data = 8'h00;
 4792 : data = 8'h00;
 4793 : data = 8'h00;
 4794 : data = 8'h00;
 4795 : data = 8'h00;
 4796 : data = 8'h00;
 4797 : data = 8'h00;
 4798 : data = 8'h00;
 4799 : data = 8'h00;
 4800 : data = 8'h00;
 4801 : data = 8'h00;
 4802 : data = 8'h00;
 4803 : data = 8'h00;
 4804 : data = 8'h00;
 4805 : data = 8'h00;
 4806 : data = 8'h00;
 4807 : data = 8'h00;
 4808 : data = 8'h00;
 4809 : data = 8'h00;
 4810 : data = 8'h00;
 4811 : data = 8'h00;
 4812 : data = 8'h00;
 4813 : data = 8'h00;
 4814 : data = 8'h00;
 4815 : data = 8'h00;
 4816 : data = 8'h00;
 4817 : data = 8'h00;
 4818 : data = 8'h00;
 4819 : data = 8'h00;
 4820 : data = 8'h00;
 4821 : data = 8'h00;
 4822 : data = 8'h00;
 4823 : data = 8'h00;
 4824 : data = 8'h00;
 4825 : data = 8'h00;
 4826 : data = 8'h00;
 4827 : data = 8'h00;
 4828 : data = 8'h00;
 4829 : data = 8'h00;
 4830 : data = 8'h00;
 4831 : data = 8'h00;
 4832 : data = 8'h00;
 4833 : data = 8'h00;
 4834 : data = 8'h00;
 4835 : data = 8'h00;
 4836 : data = 8'h00;
 4837 : data = 8'h00;
 4838 : data = 8'h00;
 4839 : data = 8'h00;
 4840 : data = 8'h00;
 4841 : data = 8'h00;
 4842 : data = 8'h00;
 4843 : data = 8'h00;
 4844 : data = 8'h00;
 4845 : data = 8'h00;
 4846 : data = 8'h00;
 4847 : data = 8'h00;
 4848 : data = 8'h00;
 4849 : data = 8'h00;
 4850 : data = 8'h00;
 4851 : data = 8'h00;
 4852 : data = 8'h00;
 4853 : data = 8'h00;
 4854 : data = 8'h00;
 4855 : data = 8'h00;
 4856 : data = 8'h00;
 4857 : data = 8'h00;
 4858 : data = 8'h00;
 4859 : data = 8'h00;
 4860 : data = 8'h00;
 4861 : data = 8'h00;
 4862 : data = 8'h00;
 4863 : data = 8'h00;
 4864 : data = 8'h00;
 4865 : data = 8'h00;
 4866 : data = 8'h00;
 4867 : data = 8'h00;
 4868 : data = 8'h00;
 4869 : data = 8'h00;
 4870 : data = 8'h00;
 4871 : data = 8'h00;
 4872 : data = 8'h00;
 4873 : data = 8'h00;
 4874 : data = 8'h00;
 4875 : data = 8'h00;
 4876 : data = 8'h00;
 4877 : data = 8'h00;
 4878 : data = 8'h00;
 4879 : data = 8'h00;
 4880 : data = 8'h00;
 4881 : data = 8'h00;
 4882 : data = 8'h00;
 4883 : data = 8'h00;
 4884 : data = 8'h00;
 4885 : data = 8'h00;
 4886 : data = 8'h00;
 4887 : data = 8'h00;
 4888 : data = 8'h00;
 4889 : data = 8'h00;
 4890 : data = 8'h00;
 4891 : data = 8'h00;
 4892 : data = 8'h00;
 4893 : data = 8'h00;
 4894 : data = 8'h00;
 4895 : data = 8'h00;
 4896 : data = 8'h00;
 4897 : data = 8'h00;
 4898 : data = 8'h00;
 4899 : data = 8'h00;
 4900 : data = 8'h00;
 4901 : data = 8'h00;
 4902 : data = 8'h00;
 4903 : data = 8'h00;
 4904 : data = 8'h00;
 4905 : data = 8'h00;
 4906 : data = 8'h00;
 4907 : data = 8'h00;
 4908 : data = 8'h00;
 4909 : data = 8'h00;
 4910 : data = 8'h00;
 4911 : data = 8'h00;
 4912 : data = 8'h00;
 4913 : data = 8'h00;
 4914 : data = 8'h00;
 4915 : data = 8'h00;
 4916 : data = 8'h00;
 4917 : data = 8'h00;
 4918 : data = 8'h00;
 4919 : data = 8'h00;
 4920 : data = 8'h00;
 4921 : data = 8'h00;
 4922 : data = 8'h00;
 4923 : data = 8'h00;
 4924 : data = 8'h00;
 4925 : data = 8'h00;
 4926 : data = 8'h00;
 4927 : data = 8'h00;
 4928 : data = 8'h00;
 4929 : data = 8'h00;
 4930 : data = 8'h00;
 4931 : data = 8'h00;
 4932 : data = 8'h00;
 4933 : data = 8'h00;
 4934 : data = 8'h00;
 4935 : data = 8'h00;
 4936 : data = 8'h00;
 4937 : data = 8'h00;
 4938 : data = 8'h00;
 4939 : data = 8'h00;
 4940 : data = 8'h00;
 4941 : data = 8'h00;
 4942 : data = 8'h00;
 4943 : data = 8'h00;
 4944 : data = 8'h00;
 4945 : data = 8'h00;
 4946 : data = 8'h00;
 4947 : data = 8'h00;
 4948 : data = 8'h00;
 4949 : data = 8'h00;
 4950 : data = 8'h00;
 4951 : data = 8'h00;
 4952 : data = 8'h00;
 4953 : data = 8'h00;
 4954 : data = 8'h00;
 4955 : data = 8'h00;
 4956 : data = 8'h00;
 4957 : data = 8'h00;
 4958 : data = 8'h00;
 4959 : data = 8'h00;
 4960 : data = 8'h00;
 4961 : data = 8'h00;
 4962 : data = 8'h00;
 4963 : data = 8'h00;
 4964 : data = 8'h00;
 4965 : data = 8'h00;
 4966 : data = 8'h00;
 4967 : data = 8'h00;
 4968 : data = 8'h00;
 4969 : data = 8'h00;
 4970 : data = 8'h00;
 4971 : data = 8'h00;
 4972 : data = 8'h00;
 4973 : data = 8'h00;
 4974 : data = 8'h00;
 4975 : data = 8'h00;
 4976 : data = 8'h00;
 4977 : data = 8'h00;
 4978 : data = 8'h00;
 4979 : data = 8'h00;
 4980 : data = 8'h00;
 4981 : data = 8'h00;
 4982 : data = 8'h00;
 4983 : data = 8'h00;
 4984 : data = 8'h00;
 4985 : data = 8'h00;
 4986 : data = 8'h00;
 4987 : data = 8'h00;
 4988 : data = 8'h00;
 4989 : data = 8'h00;
 4990 : data = 8'h00;
 4991 : data = 8'h00;
 4992 : data = 8'h00;
 4993 : data = 8'h00;
 4994 : data = 8'h00;
 4995 : data = 8'h00;
 4996 : data = 8'h00;
 4997 : data = 8'h00;
 4998 : data = 8'h00;
 4999 : data = 8'h00;
 5000 : data = 8'h00;
 5001 : data = 8'h00;
 5002 : data = 8'h00;
 5003 : data = 8'h00;
 5004 : data = 8'h00;
 5005 : data = 8'h00;
 5006 : data = 8'h00;
 5007 : data = 8'h00;
 5008 : data = 8'h00;
 5009 : data = 8'h00;
 5010 : data = 8'h00;
 5011 : data = 8'h00;
 5012 : data = 8'h00;
 5013 : data = 8'h00;
 5014 : data = 8'h00;
 5015 : data = 8'h00;
 5016 : data = 8'h00;
 5017 : data = 8'h00;
 5018 : data = 8'h00;
 5019 : data = 8'h00;
 5020 : data = 8'h00;
 5021 : data = 8'h00;
 5022 : data = 8'h00;
 5023 : data = 8'h00;
 5024 : data = 8'h00;
 5025 : data = 8'h00;
 5026 : data = 8'h00;
 5027 : data = 8'h00;
 5028 : data = 8'h00;
 5029 : data = 8'h00;
 5030 : data = 8'h00;
 5031 : data = 8'h00;
 5032 : data = 8'h00;
 5033 : data = 8'h00;
 5034 : data = 8'h00;
 5035 : data = 8'h00;
 5036 : data = 8'h00;
 5037 : data = 8'h00;
 5038 : data = 8'h00;
 5039 : data = 8'h00;
 5040 : data = 8'h00;
 5041 : data = 8'h00;
 5042 : data = 8'h00;
 5043 : data = 8'h00;
 5044 : data = 8'h00;
 5045 : data = 8'h00;
 5046 : data = 8'h00;
 5047 : data = 8'h00;
 5048 : data = 8'h00;
 5049 : data = 8'h00;
 5050 : data = 8'h00;
 5051 : data = 8'h00;
 5052 : data = 8'h00;
 5053 : data = 8'h00;
 5054 : data = 8'h00;
 5055 : data = 8'h00;
 5056 : data = 8'h00;
 5057 : data = 8'h00;
 5058 : data = 8'h00;
 5059 : data = 8'h00;
 5060 : data = 8'h00;
 5061 : data = 8'h00;
 5062 : data = 8'h00;
 5063 : data = 8'h00;
 5064 : data = 8'h00;
 5065 : data = 8'h00;
 5066 : data = 8'h00;
 5067 : data = 8'h00;
 5068 : data = 8'h00;
 5069 : data = 8'h00;
 5070 : data = 8'h00;
 5071 : data = 8'h00;
 5072 : data = 8'h00;
 5073 : data = 8'h00;
 5074 : data = 8'h00;
 5075 : data = 8'h00;
 5076 : data = 8'h00;
 5077 : data = 8'h00;
 5078 : data = 8'h00;
 5079 : data = 8'h00;
 5080 : data = 8'h00;
 5081 : data = 8'h00;
 5082 : data = 8'h00;
 5083 : data = 8'h00;
 5084 : data = 8'h00;
 5085 : data = 8'h00;
 5086 : data = 8'h00;
 5087 : data = 8'h00;
 5088 : data = 8'h00;
 5089 : data = 8'h00;
 5090 : data = 8'h00;
 5091 : data = 8'h00;
 5092 : data = 8'h00;
 5093 : data = 8'h00;
 5094 : data = 8'h00;
 5095 : data = 8'h00;
 5096 : data = 8'h00;
 5097 : data = 8'h00;
 5098 : data = 8'h00;
 5099 : data = 8'h00;
 5100 : data = 8'h00;
 5101 : data = 8'h00;
 5102 : data = 8'h00;
 5103 : data = 8'h00;
 5104 : data = 8'h00;
 5105 : data = 8'h00;
 5106 : data = 8'h00;
 5107 : data = 8'h00;
 5108 : data = 8'h00;
 5109 : data = 8'h00;
 5110 : data = 8'h00;
 5111 : data = 8'h00;
 5112 : data = 8'h00;
 5113 : data = 8'h00;
 5114 : data = 8'h00;
 5115 : data = 8'h00;
 5116 : data = 8'h00;
 5117 : data = 8'h00;
 5118 : data = 8'h00;
 5119 : data = 8'h00;
 5120 : data = 8'h00;
 5121 : data = 8'h00;
 5122 : data = 8'h00;
 5123 : data = 8'h00;
 5124 : data = 8'h00;
 5125 : data = 8'h00;
 5126 : data = 8'h00;
 5127 : data = 8'h00;
 5128 : data = 8'h00;
 5129 : data = 8'h00;
 5130 : data = 8'h00;
 5131 : data = 8'h00;
 5132 : data = 8'h00;
 5133 : data = 8'h00;
 5134 : data = 8'h00;
 5135 : data = 8'h00;
 5136 : data = 8'h00;
 5137 : data = 8'h00;
 5138 : data = 8'h00;
 5139 : data = 8'h00;
 5140 : data = 8'h00;
 5141 : data = 8'h00;
 5142 : data = 8'h00;
 5143 : data = 8'h00;
 5144 : data = 8'h00;
 5145 : data = 8'h00;
 5146 : data = 8'h00;
 5147 : data = 8'h00;
 5148 : data = 8'h00;
 5149 : data = 8'h00;
 5150 : data = 8'h00;
 5151 : data = 8'h00;
 5152 : data = 8'h00;
 5153 : data = 8'h00;
 5154 : data = 8'h00;
 5155 : data = 8'h00;
 5156 : data = 8'h00;
 5157 : data = 8'h00;
 5158 : data = 8'h00;
 5159 : data = 8'h00;
 5160 : data = 8'h00;
 5161 : data = 8'h00;
 5162 : data = 8'h00;
 5163 : data = 8'h00;
 5164 : data = 8'h00;
 5165 : data = 8'h00;
 5166 : data = 8'h00;
 5167 : data = 8'h00;
 5168 : data = 8'h00;
 5169 : data = 8'h00;
 5170 : data = 8'h00;
 5171 : data = 8'h00;
 5172 : data = 8'h00;
 5173 : data = 8'h00;
 5174 : data = 8'h00;
 5175 : data = 8'h00;
 5176 : data = 8'h00;
 5177 : data = 8'h00;
 5178 : data = 8'h00;
 5179 : data = 8'h00;
 5180 : data = 8'h00;
 5181 : data = 8'h00;
 5182 : data = 8'h00;
 5183 : data = 8'h00;
 5184 : data = 8'h00;
 5185 : data = 8'h00;
 5186 : data = 8'h00;
 5187 : data = 8'h00;
 5188 : data = 8'h00;
 5189 : data = 8'h00;
 5190 : data = 8'h00;
 5191 : data = 8'h00;
 5192 : data = 8'h00;
 5193 : data = 8'h00;
 5194 : data = 8'h00;
 5195 : data = 8'h00;
 5196 : data = 8'h00;
 5197 : data = 8'h00;
 5198 : data = 8'h00;
 5199 : data = 8'h00;
 5200 : data = 8'h00;
 5201 : data = 8'h00;
 5202 : data = 8'h00;
 5203 : data = 8'h00;
 5204 : data = 8'h00;
 5205 : data = 8'h00;
 5206 : data = 8'h00;
 5207 : data = 8'h00;
 5208 : data = 8'h00;
 5209 : data = 8'h00;
 5210 : data = 8'h00;
 5211 : data = 8'h00;
 5212 : data = 8'h00;
 5213 : data = 8'h00;
 5214 : data = 8'h00;
 5215 : data = 8'h00;
 5216 : data = 8'h00;
 5217 : data = 8'h00;
 5218 : data = 8'h00;
 5219 : data = 8'h00;
 5220 : data = 8'h00;
 5221 : data = 8'h00;
 5222 : data = 8'h00;
 5223 : data = 8'h00;
 5224 : data = 8'h00;
 5225 : data = 8'h00;
 5226 : data = 8'h00;
 5227 : data = 8'h00;
 5228 : data = 8'h00;
 5229 : data = 8'h00;
 5230 : data = 8'h00;
 5231 : data = 8'h00;
 5232 : data = 8'h00;
 5233 : data = 8'h00;
 5234 : data = 8'h00;
 5235 : data = 8'h00;
 5236 : data = 8'h00;
 5237 : data = 8'h00;
 5238 : data = 8'h00;
 5239 : data = 8'h00;
 5240 : data = 8'h00;
 5241 : data = 8'h00;
 5242 : data = 8'h00;
 5243 : data = 8'h00;
 5244 : data = 8'h00;
 5245 : data = 8'h00;
 5246 : data = 8'h00;
 5247 : data = 8'h00;
 5248 : data = 8'h00;
 5249 : data = 8'h00;
 5250 : data = 8'h00;
 5251 : data = 8'h00;
 5252 : data = 8'h00;
 5253 : data = 8'h00;
 5254 : data = 8'h00;
 5255 : data = 8'h00;
 5256 : data = 8'h00;
 5257 : data = 8'h00;
 5258 : data = 8'h00;
 5259 : data = 8'h00;
 5260 : data = 8'h00;
 5261 : data = 8'h00;
 5262 : data = 8'h00;
 5263 : data = 8'h00;
 5264 : data = 8'h00;
 5265 : data = 8'h00;
 5266 : data = 8'h00;
 5267 : data = 8'h00;
 5268 : data = 8'h00;
 5269 : data = 8'h00;
 5270 : data = 8'h00;
 5271 : data = 8'h00;
 5272 : data = 8'h00;
 5273 : data = 8'h00;
 5274 : data = 8'h00;
 5275 : data = 8'h00;
 5276 : data = 8'h00;
 5277 : data = 8'h00;
 5278 : data = 8'h00;
 5279 : data = 8'h00;
 5280 : data = 8'h00;
 5281 : data = 8'h00;
 5282 : data = 8'h00;
 5283 : data = 8'h00;
 5284 : data = 8'h00;
 5285 : data = 8'h00;
 5286 : data = 8'h00;
 5287 : data = 8'h00;
 5288 : data = 8'h00;
 5289 : data = 8'h00;
 5290 : data = 8'h00;
 5291 : data = 8'h00;
 5292 : data = 8'h00;
 5293 : data = 8'h00;
 5294 : data = 8'h00;
 5295 : data = 8'h00;
 5296 : data = 8'h00;
 5297 : data = 8'h00;
 5298 : data = 8'h00;
 5299 : data = 8'h00;
 5300 : data = 8'h00;
 5301 : data = 8'h00;
 5302 : data = 8'h00;
 5303 : data = 8'h00;
 5304 : data = 8'h00;
 5305 : data = 8'h00;
 5306 : data = 8'h00;
 5307 : data = 8'h00;
 5308 : data = 8'h00;
 5309 : data = 8'h00;
 5310 : data = 8'h00;
 5311 : data = 8'h00;
 5312 : data = 8'h00;
 5313 : data = 8'h00;
 5314 : data = 8'h00;
 5315 : data = 8'h00;
 5316 : data = 8'h00;
 5317 : data = 8'h00;
 5318 : data = 8'h00;
 5319 : data = 8'h00;
 5320 : data = 8'h00;
 5321 : data = 8'h00;
 5322 : data = 8'h00;
 5323 : data = 8'h00;
 5324 : data = 8'h00;
 5325 : data = 8'h00;
 5326 : data = 8'h00;
 5327 : data = 8'h00;
 5328 : data = 8'h00;
 5329 : data = 8'h00;
 5330 : data = 8'h00;
 5331 : data = 8'h00;
 5332 : data = 8'h00;
 5333 : data = 8'h00;
 5334 : data = 8'h00;
 5335 : data = 8'h00;
 5336 : data = 8'h00;
 5337 : data = 8'h00;
 5338 : data = 8'h00;
 5339 : data = 8'h00;
 5340 : data = 8'h00;
 5341 : data = 8'h00;
 5342 : data = 8'h00;
 5343 : data = 8'h00;
 5344 : data = 8'h00;
 5345 : data = 8'h00;
 5346 : data = 8'h00;
 5347 : data = 8'h00;
 5348 : data = 8'h00;
 5349 : data = 8'h00;
 5350 : data = 8'h00;
 5351 : data = 8'h00;
 5352 : data = 8'h00;
 5353 : data = 8'h00;
 5354 : data = 8'h00;
 5355 : data = 8'h00;
 5356 : data = 8'h00;
 5357 : data = 8'h00;
 5358 : data = 8'h00;
 5359 : data = 8'h00;
 5360 : data = 8'h00;
 5361 : data = 8'h00;
 5362 : data = 8'h00;
 5363 : data = 8'h00;
 5364 : data = 8'h00;
 5365 : data = 8'h00;
 5366 : data = 8'h00;
 5367 : data = 8'h00;
 5368 : data = 8'h00;
 5369 : data = 8'h00;
 5370 : data = 8'h00;
 5371 : data = 8'h00;
 5372 : data = 8'h00;
 5373 : data = 8'h00;
 5374 : data = 8'h00;
 5375 : data = 8'h00;
 5376 : data = 8'h00;
 5377 : data = 8'h00;
 5378 : data = 8'h00;
 5379 : data = 8'h00;
 5380 : data = 8'h00;
 5381 : data = 8'h00;
 5382 : data = 8'h00;
 5383 : data = 8'h00;
 5384 : data = 8'h00;
 5385 : data = 8'h00;
 5386 : data = 8'h00;
 5387 : data = 8'h00;
 5388 : data = 8'h00;
 5389 : data = 8'h00;
 5390 : data = 8'h00;
 5391 : data = 8'h00;
 5392 : data = 8'h00;
 5393 : data = 8'h00;
 5394 : data = 8'h00;
 5395 : data = 8'h00;
 5396 : data = 8'h00;
 5397 : data = 8'h00;
 5398 : data = 8'h00;
 5399 : data = 8'h00;
 5400 : data = 8'h00;
 5401 : data = 8'h00;
 5402 : data = 8'h00;
 5403 : data = 8'h00;
 5404 : data = 8'h00;
 5405 : data = 8'h00;
 5406 : data = 8'h00;
 5407 : data = 8'h00;
 5408 : data = 8'h00;
 5409 : data = 8'h00;
 5410 : data = 8'h00;
 5411 : data = 8'h00;
 5412 : data = 8'h00;
 5413 : data = 8'h00;
 5414 : data = 8'h00;
 5415 : data = 8'h00;
 5416 : data = 8'h00;
 5417 : data = 8'h00;
 5418 : data = 8'h00;
 5419 : data = 8'h00;
 5420 : data = 8'h00;
 5421 : data = 8'h00;
 5422 : data = 8'h00;
 5423 : data = 8'h00;
 5424 : data = 8'h00;
 5425 : data = 8'h00;
 5426 : data = 8'h00;
 5427 : data = 8'h00;
 5428 : data = 8'h00;
 5429 : data = 8'h00;
 5430 : data = 8'h00;
 5431 : data = 8'h00;
 5432 : data = 8'h00;
 5433 : data = 8'h00;
 5434 : data = 8'h00;
 5435 : data = 8'h00;
 5436 : data = 8'h00;
 5437 : data = 8'h00;
 5438 : data = 8'h00;
 5439 : data = 8'h00;
 5440 : data = 8'h00;
 5441 : data = 8'h00;
 5442 : data = 8'h00;
 5443 : data = 8'h00;
 5444 : data = 8'h00;
 5445 : data = 8'h00;
 5446 : data = 8'h00;
 5447 : data = 8'h00;
 5448 : data = 8'h00;
 5449 : data = 8'h00;
 5450 : data = 8'h00;
 5451 : data = 8'h00;
 5452 : data = 8'h00;
 5453 : data = 8'h00;
 5454 : data = 8'h00;
 5455 : data = 8'h00;
 5456 : data = 8'h00;
 5457 : data = 8'h00;
 5458 : data = 8'h00;
 5459 : data = 8'h00;
 5460 : data = 8'h00;
 5461 : data = 8'h00;
 5462 : data = 8'h00;
 5463 : data = 8'h00;
 5464 : data = 8'h00;
 5465 : data = 8'h00;
 5466 : data = 8'h00;
 5467 : data = 8'h00;
 5468 : data = 8'h00;
 5469 : data = 8'h00;
 5470 : data = 8'h00;
 5471 : data = 8'h00;
 5472 : data = 8'h00;
 5473 : data = 8'h00;
 5474 : data = 8'h00;
 5475 : data = 8'h00;
 5476 : data = 8'h00;
 5477 : data = 8'h00;
 5478 : data = 8'h00;
 5479 : data = 8'h00;
 5480 : data = 8'h00;
 5481 : data = 8'h00;
 5482 : data = 8'h00;
 5483 : data = 8'h00;
 5484 : data = 8'h00;
 5485 : data = 8'h00;
 5486 : data = 8'h00;
 5487 : data = 8'h00;
 5488 : data = 8'h00;
 5489 : data = 8'h00;
 5490 : data = 8'h00;
 5491 : data = 8'h00;
 5492 : data = 8'h00;
 5493 : data = 8'h00;
 5494 : data = 8'h00;
 5495 : data = 8'h00;
 5496 : data = 8'h00;
 5497 : data = 8'h00;
 5498 : data = 8'h00;
 5499 : data = 8'h00;
 5500 : data = 8'h00;
 5501 : data = 8'h00;
 5502 : data = 8'h00;
 5503 : data = 8'h00;
 5504 : data = 8'h00;
 5505 : data = 8'h00;
 5506 : data = 8'h00;
 5507 : data = 8'h00;
 5508 : data = 8'h00;
 5509 : data = 8'h00;
 5510 : data = 8'h00;
 5511 : data = 8'h00;
 5512 : data = 8'h00;
 5513 : data = 8'h00;
 5514 : data = 8'h00;
 5515 : data = 8'h00;
 5516 : data = 8'h00;
 5517 : data = 8'h00;
 5518 : data = 8'h00;
 5519 : data = 8'h00;
 5520 : data = 8'h00;
 5521 : data = 8'h00;
 5522 : data = 8'h00;
 5523 : data = 8'h00;
 5524 : data = 8'h00;
 5525 : data = 8'h00;
 5526 : data = 8'h00;
 5527 : data = 8'h00;
 5528 : data = 8'h00;
 5529 : data = 8'h00;
 5530 : data = 8'h00;
 5531 : data = 8'h00;
 5532 : data = 8'h00;
 5533 : data = 8'h00;
 5534 : data = 8'h00;
 5535 : data = 8'h00;
 5536 : data = 8'h00;
 5537 : data = 8'h00;
 5538 : data = 8'h00;
 5539 : data = 8'h00;
 5540 : data = 8'h00;
 5541 : data = 8'h00;
 5542 : data = 8'h00;
 5543 : data = 8'h00;
 5544 : data = 8'h00;
 5545 : data = 8'h00;
 5546 : data = 8'h00;
 5547 : data = 8'h00;
 5548 : data = 8'h00;
 5549 : data = 8'h00;
 5550 : data = 8'h00;
 5551 : data = 8'h00;
 5552 : data = 8'h00;
 5553 : data = 8'h00;
 5554 : data = 8'h00;
 5555 : data = 8'h00;
 5556 : data = 8'h00;
 5557 : data = 8'h00;
 5558 : data = 8'h00;
 5559 : data = 8'h00;
 5560 : data = 8'h00;
 5561 : data = 8'h00;
 5562 : data = 8'h00;
 5563 : data = 8'h00;
 5564 : data = 8'h00;
 5565 : data = 8'h00;
 5566 : data = 8'h00;
 5567 : data = 8'h00;
 5568 : data = 8'h00;
 5569 : data = 8'h00;
 5570 : data = 8'h00;
 5571 : data = 8'h00;
 5572 : data = 8'h00;
 5573 : data = 8'h00;
 5574 : data = 8'h00;
 5575 : data = 8'h00;
 5576 : data = 8'h00;
 5577 : data = 8'h00;
 5578 : data = 8'h00;
 5579 : data = 8'h00;
 5580 : data = 8'h00;
 5581 : data = 8'h00;
 5582 : data = 8'h00;
 5583 : data = 8'h00;
 5584 : data = 8'h00;
 5585 : data = 8'h00;
 5586 : data = 8'h00;
 5587 : data = 8'h00;
 5588 : data = 8'h00;
 5589 : data = 8'h00;
 5590 : data = 8'h00;
 5591 : data = 8'h00;
 5592 : data = 8'h00;
 5593 : data = 8'h00;
 5594 : data = 8'h00;
 5595 : data = 8'h00;
 5596 : data = 8'h00;
 5597 : data = 8'h00;
 5598 : data = 8'h00;
 5599 : data = 8'h00;
 5600 : data = 8'h00;
 5601 : data = 8'h00;
 5602 : data = 8'h00;
 5603 : data = 8'h00;
 5604 : data = 8'h00;
 5605 : data = 8'h00;
 5606 : data = 8'h00;
 5607 : data = 8'h00;
 5608 : data = 8'h00;
 5609 : data = 8'h00;
 5610 : data = 8'h00;
 5611 : data = 8'h00;
 5612 : data = 8'h00;
 5613 : data = 8'h00;
 5614 : data = 8'h00;
 5615 : data = 8'h00;
 5616 : data = 8'h00;
 5617 : data = 8'h00;
 5618 : data = 8'h00;
 5619 : data = 8'h00;
 5620 : data = 8'h00;
 5621 : data = 8'h00;
 5622 : data = 8'h00;
 5623 : data = 8'h00;
 5624 : data = 8'h00;
 5625 : data = 8'h00;
 5626 : data = 8'h00;
 5627 : data = 8'h00;
 5628 : data = 8'h00;
 5629 : data = 8'h00;
 5630 : data = 8'h00;
 5631 : data = 8'h00;
 5632 : data = 8'h00;
 5633 : data = 8'h00;
 5634 : data = 8'h00;
 5635 : data = 8'h00;
 5636 : data = 8'h00;
 5637 : data = 8'h00;
 5638 : data = 8'h00;
 5639 : data = 8'h00;
 5640 : data = 8'h00;
 5641 : data = 8'h00;
 5642 : data = 8'h00;
 5643 : data = 8'h00;
 5644 : data = 8'h00;
 5645 : data = 8'h00;
 5646 : data = 8'h00;
 5647 : data = 8'h00;
 5648 : data = 8'h00;
 5649 : data = 8'h00;
 5650 : data = 8'h00;
 5651 : data = 8'h00;
 5652 : data = 8'h00;
 5653 : data = 8'h00;
 5654 : data = 8'h00;
 5655 : data = 8'h00;
 5656 : data = 8'h00;
 5657 : data = 8'h00;
 5658 : data = 8'h00;
 5659 : data = 8'h00;
 5660 : data = 8'h00;
 5661 : data = 8'h00;
 5662 : data = 8'h00;
 5663 : data = 8'h00;
 5664 : data = 8'h00;
 5665 : data = 8'h00;
 5666 : data = 8'h00;
 5667 : data = 8'h00;
 5668 : data = 8'h00;
 5669 : data = 8'h00;
 5670 : data = 8'h00;
 5671 : data = 8'h00;
 5672 : data = 8'h00;
 5673 : data = 8'h00;
 5674 : data = 8'h00;
 5675 : data = 8'h00;
 5676 : data = 8'h00;
 5677 : data = 8'h00;
 5678 : data = 8'h00;
 5679 : data = 8'h00;
 5680 : data = 8'h00;
 5681 : data = 8'h00;
 5682 : data = 8'h00;
 5683 : data = 8'h00;
 5684 : data = 8'h00;
 5685 : data = 8'h00;
 5686 : data = 8'h00;
 5687 : data = 8'h00;
 5688 : data = 8'h00;
 5689 : data = 8'h00;
 5690 : data = 8'h00;
 5691 : data = 8'h00;
 5692 : data = 8'h00;
 5693 : data = 8'h00;
 5694 : data = 8'h00;
 5695 : data = 8'h00;
 5696 : data = 8'h00;
 5697 : data = 8'h00;
 5698 : data = 8'h00;
 5699 : data = 8'h00;
 5700 : data = 8'h00;
 5701 : data = 8'h00;
 5702 : data = 8'h00;
 5703 : data = 8'h00;
 5704 : data = 8'h00;
 5705 : data = 8'h00;
 5706 : data = 8'h00;
 5707 : data = 8'h00;
 5708 : data = 8'h00;
 5709 : data = 8'h00;
 5710 : data = 8'h00;
 5711 : data = 8'h00;
 5712 : data = 8'h00;
 5713 : data = 8'h00;
 5714 : data = 8'h00;
 5715 : data = 8'h00;
 5716 : data = 8'h00;
 5717 : data = 8'h00;
 5718 : data = 8'h00;
 5719 : data = 8'h00;
 5720 : data = 8'h00;
 5721 : data = 8'h00;
 5722 : data = 8'h00;
 5723 : data = 8'h00;
 5724 : data = 8'h00;
 5725 : data = 8'h00;
 5726 : data = 8'h00;
 5727 : data = 8'h00;
 5728 : data = 8'h00;
 5729 : data = 8'h00;
 5730 : data = 8'h00;
 5731 : data = 8'h00;
 5732 : data = 8'h00;
 5733 : data = 8'h00;
 5734 : data = 8'h00;
 5735 : data = 8'h00;
 5736 : data = 8'h00;
 5737 : data = 8'h00;
 5738 : data = 8'h00;
 5739 : data = 8'h00;
 5740 : data = 8'h00;
 5741 : data = 8'h00;
 5742 : data = 8'h00;
 5743 : data = 8'h00;
 5744 : data = 8'h00;
 5745 : data = 8'h00;
 5746 : data = 8'h00;
 5747 : data = 8'h00;
 5748 : data = 8'h00;
 5749 : data = 8'h00;
 5750 : data = 8'h00;
 5751 : data = 8'h00;
 5752 : data = 8'h00;
 5753 : data = 8'h00;
 5754 : data = 8'h00;
 5755 : data = 8'h00;
 5756 : data = 8'h00;
 5757 : data = 8'h00;
 5758 : data = 8'h00;
 5759 : data = 8'h00;
 5760 : data = 8'h00;
 5761 : data = 8'h00;
 5762 : data = 8'h00;
 5763 : data = 8'h00;
 5764 : data = 8'h00;
 5765 : data = 8'h00;
 5766 : data = 8'h00;
 5767 : data = 8'h00;
 5768 : data = 8'h00;
 5769 : data = 8'h00;
 5770 : data = 8'h00;
 5771 : data = 8'h00;
 5772 : data = 8'h00;
 5773 : data = 8'h00;
 5774 : data = 8'h00;
 5775 : data = 8'h00;
 5776 : data = 8'h00;
 5777 : data = 8'h00;
 5778 : data = 8'h00;
 5779 : data = 8'h00;
 5780 : data = 8'h00;
 5781 : data = 8'h00;
 5782 : data = 8'h00;
 5783 : data = 8'h00;
 5784 : data = 8'h00;
 5785 : data = 8'h00;
 5786 : data = 8'h00;
 5787 : data = 8'h00;
 5788 : data = 8'h00;
 5789 : data = 8'h00;
 5790 : data = 8'h00;
 5791 : data = 8'h00;
 5792 : data = 8'h00;
 5793 : data = 8'h00;
 5794 : data = 8'h00;
 5795 : data = 8'h00;
 5796 : data = 8'h00;
 5797 : data = 8'h00;
 5798 : data = 8'h00;
 5799 : data = 8'h00;
 5800 : data = 8'h00;
 5801 : data = 8'h00;
 5802 : data = 8'h00;
 5803 : data = 8'h00;
 5804 : data = 8'h00;
 5805 : data = 8'h00;
 5806 : data = 8'h00;
 5807 : data = 8'h00;
 5808 : data = 8'h00;
 5809 : data = 8'h00;
 5810 : data = 8'h00;
 5811 : data = 8'h00;
 5812 : data = 8'h00;
 5813 : data = 8'h00;
 5814 : data = 8'h00;
 5815 : data = 8'h00;
 5816 : data = 8'h00;
 5817 : data = 8'h00;
 5818 : data = 8'h00;
 5819 : data = 8'h00;
 5820 : data = 8'h00;
 5821 : data = 8'h00;
 5822 : data = 8'h00;
 5823 : data = 8'h00;
 5824 : data = 8'h00;
 5825 : data = 8'h00;
 5826 : data = 8'h00;
 5827 : data = 8'h00;
 5828 : data = 8'h00;
 5829 : data = 8'h00;
 5830 : data = 8'h00;
 5831 : data = 8'h00;
 5832 : data = 8'h00;
 5833 : data = 8'h00;
 5834 : data = 8'h00;
 5835 : data = 8'h00;
 5836 : data = 8'h00;
 5837 : data = 8'h00;
 5838 : data = 8'h00;
 5839 : data = 8'h00;
 5840 : data = 8'h00;
 5841 : data = 8'h00;
 5842 : data = 8'h00;
 5843 : data = 8'h00;
 5844 : data = 8'h00;
 5845 : data = 8'h00;
 5846 : data = 8'h00;
 5847 : data = 8'h00;
 5848 : data = 8'h00;
 5849 : data = 8'h00;
 5850 : data = 8'h00;
 5851 : data = 8'h00;
 5852 : data = 8'h00;
 5853 : data = 8'h00;
 5854 : data = 8'h00;
 5855 : data = 8'h00;
 5856 : data = 8'h00;
 5857 : data = 8'h00;
 5858 : data = 8'h00;
 5859 : data = 8'h00;
 5860 : data = 8'h00;
 5861 : data = 8'h00;
 5862 : data = 8'h00;
 5863 : data = 8'h00;
 5864 : data = 8'h00;
 5865 : data = 8'h00;
 5866 : data = 8'h00;
 5867 : data = 8'h00;
 5868 : data = 8'h00;
 5869 : data = 8'h00;
 5870 : data = 8'h00;
 5871 : data = 8'h00;
 5872 : data = 8'h00;
 5873 : data = 8'h00;
 5874 : data = 8'h00;
 5875 : data = 8'h00;
 5876 : data = 8'h00;
 5877 : data = 8'h00;
 5878 : data = 8'h00;
 5879 : data = 8'h00;
 5880 : data = 8'h00;
 5881 : data = 8'h00;
 5882 : data = 8'h00;
 5883 : data = 8'h00;
 5884 : data = 8'h00;
 5885 : data = 8'h00;
 5886 : data = 8'h00;
 5887 : data = 8'h00;
 5888 : data = 8'h00;
 5889 : data = 8'h00;
 5890 : data = 8'h00;
 5891 : data = 8'h00;
 5892 : data = 8'h00;
 5893 : data = 8'h00;
 5894 : data = 8'h00;
 5895 : data = 8'h00;
 5896 : data = 8'h00;
 5897 : data = 8'h00;
 5898 : data = 8'h00;
 5899 : data = 8'h00;
 5900 : data = 8'h00;
 5901 : data = 8'h00;
 5902 : data = 8'h00;
 5903 : data = 8'h00;
 5904 : data = 8'h00;
 5905 : data = 8'h00;
 5906 : data = 8'h00;
 5907 : data = 8'h00;
 5908 : data = 8'h00;
 5909 : data = 8'h00;
 5910 : data = 8'h00;
 5911 : data = 8'h00;
 5912 : data = 8'h00;
 5913 : data = 8'h00;
 5914 : data = 8'h00;
 5915 : data = 8'h00;
 5916 : data = 8'h00;
 5917 : data = 8'h00;
 5918 : data = 8'h00;
 5919 : data = 8'h00;
 5920 : data = 8'h00;
 5921 : data = 8'h00;
 5922 : data = 8'h00;
 5923 : data = 8'h00;
 5924 : data = 8'h00;
 5925 : data = 8'h00;
 5926 : data = 8'h00;
 5927 : data = 8'h00;
 5928 : data = 8'h00;
 5929 : data = 8'h00;
 5930 : data = 8'h00;
 5931 : data = 8'h00;
 5932 : data = 8'h00;
 5933 : data = 8'h00;
 5934 : data = 8'h00;
 5935 : data = 8'h00;
 5936 : data = 8'h00;
 5937 : data = 8'h00;
 5938 : data = 8'h00;
 5939 : data = 8'h00;
 5940 : data = 8'h00;
 5941 : data = 8'h00;
 5942 : data = 8'h00;
 5943 : data = 8'h00;
 5944 : data = 8'h00;
 5945 : data = 8'h00;
 5946 : data = 8'h00;
 5947 : data = 8'h00;
 5948 : data = 8'h00;
 5949 : data = 8'h00;
 5950 : data = 8'h00;
 5951 : data = 8'h00;
 5952 : data = 8'h00;
 5953 : data = 8'h00;
 5954 : data = 8'h00;
 5955 : data = 8'h00;
 5956 : data = 8'h00;
 5957 : data = 8'h00;
 5958 : data = 8'h00;
 5959 : data = 8'h00;
 5960 : data = 8'h00;
 5961 : data = 8'h00;
 5962 : data = 8'h00;
 5963 : data = 8'h00;
 5964 : data = 8'h00;
 5965 : data = 8'h00;
 5966 : data = 8'h00;
 5967 : data = 8'h00;
 5968 : data = 8'h00;
 5969 : data = 8'h00;
 5970 : data = 8'h00;
 5971 : data = 8'h00;
 5972 : data = 8'h00;
 5973 : data = 8'h00;
 5974 : data = 8'h00;
 5975 : data = 8'h00;
 5976 : data = 8'h00;
 5977 : data = 8'h00;
 5978 : data = 8'h00;
 5979 : data = 8'h00;
 5980 : data = 8'h00;
 5981 : data = 8'h00;
 5982 : data = 8'h00;
 5983 : data = 8'h00;
 5984 : data = 8'h00;
 5985 : data = 8'h00;
 5986 : data = 8'h00;
 5987 : data = 8'h00;
 5988 : data = 8'h00;
 5989 : data = 8'h00;
 5990 : data = 8'h00;
 5991 : data = 8'h00;
 5992 : data = 8'h00;
 5993 : data = 8'h00;
 5994 : data = 8'h00;
 5995 : data = 8'h00;
 5996 : data = 8'h00;
 5997 : data = 8'h00;
 5998 : data = 8'h00;
 5999 : data = 8'h00;
 6000 : data = 8'h00;
 6001 : data = 8'h00;
 6002 : data = 8'h00;
 6003 : data = 8'h00;
 6004 : data = 8'h00;
 6005 : data = 8'h00;
 6006 : data = 8'h00;
 6007 : data = 8'h00;
 6008 : data = 8'h00;
 6009 : data = 8'h00;
 6010 : data = 8'h00;
 6011 : data = 8'h00;
 6012 : data = 8'h00;
 6013 : data = 8'h00;
 6014 : data = 8'h00;
 6015 : data = 8'h00;
 6016 : data = 8'h00;
 6017 : data = 8'h00;
 6018 : data = 8'h00;
 6019 : data = 8'h00;
 6020 : data = 8'h00;
 6021 : data = 8'h00;
 6022 : data = 8'h00;
 6023 : data = 8'h00;
 6024 : data = 8'h00;
 6025 : data = 8'h00;
 6026 : data = 8'h00;
 6027 : data = 8'h00;
 6028 : data = 8'h00;
 6029 : data = 8'h00;
 6030 : data = 8'h00;
 6031 : data = 8'h00;
 6032 : data = 8'h00;
 6033 : data = 8'h00;
 6034 : data = 8'h00;
 6035 : data = 8'h00;
 6036 : data = 8'h00;
 6037 : data = 8'h00;
 6038 : data = 8'h00;
 6039 : data = 8'h00;
 6040 : data = 8'h00;
 6041 : data = 8'h00;
 6042 : data = 8'h00;
 6043 : data = 8'h00;
 6044 : data = 8'h00;
 6045 : data = 8'h00;
 6046 : data = 8'h00;
 6047 : data = 8'h00;
 6048 : data = 8'h00;
 6049 : data = 8'h00;
 6050 : data = 8'h00;
 6051 : data = 8'h00;
 6052 : data = 8'h00;
 6053 : data = 8'h00;
 6054 : data = 8'h00;
 6055 : data = 8'h00;
 6056 : data = 8'h00;
 6057 : data = 8'h00;
 6058 : data = 8'h00;
 6059 : data = 8'h00;
 6060 : data = 8'h00;
 6061 : data = 8'h00;
 6062 : data = 8'h00;
 6063 : data = 8'h00;
 6064 : data = 8'h00;
 6065 : data = 8'h00;
 6066 : data = 8'h00;
 6067 : data = 8'h00;
 6068 : data = 8'h00;
 6069 : data = 8'h00;
 6070 : data = 8'h00;
 6071 : data = 8'h00;
 6072 : data = 8'h00;
 6073 : data = 8'h00;
 6074 : data = 8'h00;
 6075 : data = 8'h00;
 6076 : data = 8'h00;
 6077 : data = 8'h00;
 6078 : data = 8'h00;
 6079 : data = 8'h00;
 6080 : data = 8'h00;
 6081 : data = 8'h00;
 6082 : data = 8'h00;
 6083 : data = 8'h00;
 6084 : data = 8'h00;
 6085 : data = 8'h00;
 6086 : data = 8'h00;
 6087 : data = 8'h00;
 6088 : data = 8'h00;
 6089 : data = 8'h00;
 6090 : data = 8'h00;
 6091 : data = 8'h00;
 6092 : data = 8'h00;
 6093 : data = 8'h00;
 6094 : data = 8'h00;
 6095 : data = 8'h00;
 6096 : data = 8'h00;
 6097 : data = 8'h00;
 6098 : data = 8'h00;
 6099 : data = 8'h00;
 6100 : data = 8'h00;
 6101 : data = 8'h00;
 6102 : data = 8'h00;
 6103 : data = 8'h00;
 6104 : data = 8'h00;
 6105 : data = 8'h00;
 6106 : data = 8'h00;
 6107 : data = 8'h00;
 6108 : data = 8'h00;
 6109 : data = 8'h00;
 6110 : data = 8'h00;
 6111 : data = 8'h00;
 6112 : data = 8'h00;
 6113 : data = 8'h00;
 6114 : data = 8'h00;
 6115 : data = 8'h00;
 6116 : data = 8'h00;
 6117 : data = 8'h00;
 6118 : data = 8'h00;
 6119 : data = 8'h00;
 6120 : data = 8'h00;
 6121 : data = 8'h00;
 6122 : data = 8'h00;
 6123 : data = 8'h00;
 6124 : data = 8'h00;
 6125 : data = 8'h00;
 6126 : data = 8'h00;
 6127 : data = 8'h00;
 6128 : data = 8'h00;
 6129 : data = 8'h00;
 6130 : data = 8'h00;
 6131 : data = 8'h00;
 6132 : data = 8'h00;
 6133 : data = 8'h00;
 6134 : data = 8'h00;
 6135 : data = 8'h00;
 6136 : data = 8'h00;
 6137 : data = 8'h00;
 6138 : data = 8'h00;
 6139 : data = 8'h00;
 6140 : data = 8'h00;
 6141 : data = 8'h00;
 6142 : data = 8'h00;
 6143 : data = 8'h00;
 6144 : data = 8'h00;
 6145 : data = 8'h00;
 6146 : data = 8'h00;
 6147 : data = 8'h00;
 6148 : data = 8'h00;
 6149 : data = 8'h00;
 6150 : data = 8'h00;
 6151 : data = 8'h00;
 6152 : data = 8'h00;
 6153 : data = 8'h00;
 6154 : data = 8'h00;
 6155 : data = 8'h00;
 6156 : data = 8'h00;
 6157 : data = 8'h00;
 6158 : data = 8'h00;
 6159 : data = 8'h00;
 6160 : data = 8'h00;
 6161 : data = 8'h00;
 6162 : data = 8'h00;
 6163 : data = 8'h00;
 6164 : data = 8'h00;
 6165 : data = 8'h00;
 6166 : data = 8'h00;
 6167 : data = 8'h00;
 6168 : data = 8'h00;
 6169 : data = 8'h00;
 6170 : data = 8'h00;
 6171 : data = 8'h00;
 6172 : data = 8'h00;
 6173 : data = 8'h00;
 6174 : data = 8'h00;
 6175 : data = 8'h00;
 6176 : data = 8'h00;
 6177 : data = 8'h00;
 6178 : data = 8'h00;
 6179 : data = 8'h00;
 6180 : data = 8'h00;
 6181 : data = 8'h00;
 6182 : data = 8'h00;
 6183 : data = 8'h00;
 6184 : data = 8'h00;
 6185 : data = 8'h00;
 6186 : data = 8'h00;
 6187 : data = 8'h00;
 6188 : data = 8'h00;
 6189 : data = 8'h00;
 6190 : data = 8'h00;
 6191 : data = 8'h00;
 6192 : data = 8'h00;
 6193 : data = 8'h00;
 6194 : data = 8'h00;
 6195 : data = 8'h00;
 6196 : data = 8'h00;
 6197 : data = 8'h00;
 6198 : data = 8'h00;
 6199 : data = 8'h00;
 6200 : data = 8'h00;
 6201 : data = 8'h00;
 6202 : data = 8'h00;
 6203 : data = 8'h00;
 6204 : data = 8'h00;
 6205 : data = 8'h00;
 6206 : data = 8'h00;
 6207 : data = 8'h00;
 6208 : data = 8'h00;
 6209 : data = 8'h00;
 6210 : data = 8'h00;
 6211 : data = 8'h00;
 6212 : data = 8'h00;
 6213 : data = 8'h00;
 6214 : data = 8'h00;
 6215 : data = 8'h00;
 6216 : data = 8'h00;
 6217 : data = 8'h00;
 6218 : data = 8'h00;
 6219 : data = 8'h00;
 6220 : data = 8'h00;
 6221 : data = 8'h00;
 6222 : data = 8'h00;
 6223 : data = 8'h00;
 6224 : data = 8'h00;
 6225 : data = 8'h00;
 6226 : data = 8'h00;
 6227 : data = 8'h00;
 6228 : data = 8'h00;
 6229 : data = 8'h00;
 6230 : data = 8'h00;
 6231 : data = 8'h00;
 6232 : data = 8'h00;
 6233 : data = 8'h00;
 6234 : data = 8'h00;
 6235 : data = 8'h00;
 6236 : data = 8'h00;
 6237 : data = 8'h00;
 6238 : data = 8'h00;
 6239 : data = 8'h00;
 6240 : data = 8'h00;
 6241 : data = 8'h00;
 6242 : data = 8'h00;
 6243 : data = 8'h00;
 6244 : data = 8'h00;
 6245 : data = 8'h00;
 6246 : data = 8'h00;
 6247 : data = 8'h00;
 6248 : data = 8'h00;
 6249 : data = 8'h00;
 6250 : data = 8'h00;
 6251 : data = 8'h00;
 6252 : data = 8'h00;
 6253 : data = 8'h00;
 6254 : data = 8'h00;
 6255 : data = 8'h00;
 6256 : data = 8'h00;
 6257 : data = 8'h00;
 6258 : data = 8'h00;
 6259 : data = 8'h00;
 6260 : data = 8'h00;
 6261 : data = 8'h00;
 6262 : data = 8'h00;
 6263 : data = 8'h00;
 6264 : data = 8'h00;
 6265 : data = 8'h00;
 6266 : data = 8'h00;
 6267 : data = 8'h00;
 6268 : data = 8'h00;
 6269 : data = 8'h00;
 6270 : data = 8'h00;
 6271 : data = 8'h00;
 6272 : data = 8'h00;
 6273 : data = 8'h00;
 6274 : data = 8'h00;
 6275 : data = 8'h00;
 6276 : data = 8'h00;
 6277 : data = 8'h00;
 6278 : data = 8'h00;
 6279 : data = 8'h00;
 6280 : data = 8'h00;
 6281 : data = 8'h00;
 6282 : data = 8'h00;
 6283 : data = 8'h00;
 6284 : data = 8'h00;
 6285 : data = 8'h00;
 6286 : data = 8'h00;
 6287 : data = 8'h00;
 6288 : data = 8'h00;
 6289 : data = 8'h00;
 6290 : data = 8'h00;
 6291 : data = 8'h00;
 6292 : data = 8'h00;
 6293 : data = 8'h00;
 6294 : data = 8'h00;
 6295 : data = 8'h00;
 6296 : data = 8'h00;
 6297 : data = 8'h00;
 6298 : data = 8'h00;
 6299 : data = 8'h00;
 6300 : data = 8'h00;
 6301 : data = 8'h00;
 6302 : data = 8'h00;
 6303 : data = 8'h00;
 6304 : data = 8'h00;
 6305 : data = 8'h00;
 6306 : data = 8'h00;
 6307 : data = 8'h00;
 6308 : data = 8'h00;
 6309 : data = 8'h00;
 6310 : data = 8'h00;
 6311 : data = 8'h00;
 6312 : data = 8'h00;
 6313 : data = 8'h00;
 6314 : data = 8'h00;
 6315 : data = 8'h00;
 6316 : data = 8'h00;
 6317 : data = 8'h00;
 6318 : data = 8'h00;
 6319 : data = 8'h00;
 6320 : data = 8'h00;
 6321 : data = 8'h00;
 6322 : data = 8'h00;
 6323 : data = 8'h00;
 6324 : data = 8'h00;
 6325 : data = 8'h00;
 6326 : data = 8'h00;
 6327 : data = 8'h00;
 6328 : data = 8'h00;
 6329 : data = 8'h00;
 6330 : data = 8'h00;
 6331 : data = 8'h00;
 6332 : data = 8'h00;
 6333 : data = 8'h00;
 6334 : data = 8'h00;
 6335 : data = 8'h00;
 6336 : data = 8'h00;
 6337 : data = 8'h00;
 6338 : data = 8'h00;
 6339 : data = 8'h00;
 6340 : data = 8'h00;
 6341 : data = 8'h00;
 6342 : data = 8'h00;
 6343 : data = 8'h00;
 6344 : data = 8'h00;
 6345 : data = 8'h00;
 6346 : data = 8'h00;
 6347 : data = 8'h00;
 6348 : data = 8'h00;
 6349 : data = 8'h00;
 6350 : data = 8'h00;
 6351 : data = 8'h00;
 6352 : data = 8'h00;
 6353 : data = 8'h00;
 6354 : data = 8'h00;
 6355 : data = 8'h00;
 6356 : data = 8'h00;
 6357 : data = 8'h00;
 6358 : data = 8'h00;
 6359 : data = 8'h00;
 6360 : data = 8'h00;
 6361 : data = 8'h00;
 6362 : data = 8'h00;
 6363 : data = 8'h00;
 6364 : data = 8'h00;
 6365 : data = 8'h00;
 6366 : data = 8'h00;
 6367 : data = 8'h00;
 6368 : data = 8'h00;
 6369 : data = 8'h00;
 6370 : data = 8'h00;
 6371 : data = 8'h00;
 6372 : data = 8'h00;
 6373 : data = 8'h00;
 6374 : data = 8'h00;
 6375 : data = 8'h00;
 6376 : data = 8'h00;
 6377 : data = 8'h00;
 6378 : data = 8'h00;
 6379 : data = 8'h00;
 6380 : data = 8'h00;
 6381 : data = 8'h00;
 6382 : data = 8'h00;
 6383 : data = 8'h00;
 6384 : data = 8'h00;
 6385 : data = 8'h00;
 6386 : data = 8'h00;
 6387 : data = 8'h00;
 6388 : data = 8'h00;
 6389 : data = 8'h00;
 6390 : data = 8'h00;
 6391 : data = 8'h00;
 6392 : data = 8'h00;
 6393 : data = 8'h00;
 6394 : data = 8'h00;
 6395 : data = 8'h00;
 6396 : data = 8'h00;
 6397 : data = 8'h00;
 6398 : data = 8'h00;
 6399 : data = 8'h00;
 6400 : data = 8'h00;
 6401 : data = 8'h00;
 6402 : data = 8'h00;
 6403 : data = 8'h00;
 6404 : data = 8'h00;
 6405 : data = 8'h00;
 6406 : data = 8'h00;
 6407 : data = 8'h00;
 6408 : data = 8'h00;
 6409 : data = 8'h00;
 6410 : data = 8'h00;
 6411 : data = 8'h00;
 6412 : data = 8'h00;
 6413 : data = 8'h00;
 6414 : data = 8'h00;
 6415 : data = 8'h00;
 6416 : data = 8'h00;
 6417 : data = 8'h00;
 6418 : data = 8'h00;
 6419 : data = 8'h00;
 6420 : data = 8'h00;
 6421 : data = 8'h00;
 6422 : data = 8'h00;
 6423 : data = 8'h00;
 6424 : data = 8'h00;
 6425 : data = 8'h00;
 6426 : data = 8'h00;
 6427 : data = 8'h00;
 6428 : data = 8'h00;
 6429 : data = 8'h00;
 6430 : data = 8'h00;
 6431 : data = 8'h00;
 6432 : data = 8'h00;
 6433 : data = 8'h00;
 6434 : data = 8'h00;
 6435 : data = 8'h00;
 6436 : data = 8'h00;
 6437 : data = 8'h00;
 6438 : data = 8'h00;
 6439 : data = 8'h00;
 6440 : data = 8'h00;
 6441 : data = 8'h00;
 6442 : data = 8'h00;
 6443 : data = 8'h00;
 6444 : data = 8'h00;
 6445 : data = 8'h00;
 6446 : data = 8'h00;
 6447 : data = 8'h00;
 6448 : data = 8'h00;
 6449 : data = 8'h00;
 6450 : data = 8'h00;
 6451 : data = 8'h00;
 6452 : data = 8'h00;
 6453 : data = 8'h00;
 6454 : data = 8'h00;
 6455 : data = 8'h00;
 6456 : data = 8'h00;
 6457 : data = 8'h00;
 6458 : data = 8'h00;
 6459 : data = 8'h00;
 6460 : data = 8'h00;
 6461 : data = 8'h00;
 6462 : data = 8'h00;
 6463 : data = 8'h00;
 6464 : data = 8'h00;
 6465 : data = 8'h00;
 6466 : data = 8'h00;
 6467 : data = 8'h00;
 6468 : data = 8'h00;
 6469 : data = 8'h00;
 6470 : data = 8'h00;
 6471 : data = 8'h00;
 6472 : data = 8'h00;
 6473 : data = 8'h00;
 6474 : data = 8'h00;
 6475 : data = 8'h00;
 6476 : data = 8'h00;
 6477 : data = 8'h00;
 6478 : data = 8'h00;
 6479 : data = 8'h00;
 6480 : data = 8'h00;
 6481 : data = 8'h00;
 6482 : data = 8'h00;
 6483 : data = 8'h00;
 6484 : data = 8'h00;
 6485 : data = 8'h00;
 6486 : data = 8'h00;
 6487 : data = 8'h00;
 6488 : data = 8'h00;
 6489 : data = 8'h00;
 6490 : data = 8'h00;
 6491 : data = 8'h00;
 6492 : data = 8'h00;
 6493 : data = 8'h00;
 6494 : data = 8'h00;
 6495 : data = 8'h00;
 6496 : data = 8'h00;
 6497 : data = 8'h00;
 6498 : data = 8'h00;
 6499 : data = 8'h00;
 6500 : data = 8'h00;
 6501 : data = 8'h00;
 6502 : data = 8'h00;
 6503 : data = 8'h00;
 6504 : data = 8'h00;
 6505 : data = 8'h00;
 6506 : data = 8'h00;
 6507 : data = 8'h00;
 6508 : data = 8'h00;
 6509 : data = 8'h00;
 6510 : data = 8'h00;
 6511 : data = 8'h00;
 6512 : data = 8'h00;
 6513 : data = 8'h00;
 6514 : data = 8'h00;
 6515 : data = 8'h00;
 6516 : data = 8'h00;
 6517 : data = 8'h00;
 6518 : data = 8'h00;
 6519 : data = 8'h00;
 6520 : data = 8'h00;
 6521 : data = 8'h00;
 6522 : data = 8'h00;
 6523 : data = 8'h00;
 6524 : data = 8'h00;
 6525 : data = 8'h00;
 6526 : data = 8'h00;
 6527 : data = 8'h00;
 6528 : data = 8'h00;
 6529 : data = 8'h00;
 6530 : data = 8'h00;
 6531 : data = 8'h00;
 6532 : data = 8'h00;
 6533 : data = 8'h00;
 6534 : data = 8'h00;
 6535 : data = 8'h00;
 6536 : data = 8'h00;
 6537 : data = 8'h00;
 6538 : data = 8'h00;
 6539 : data = 8'h00;
 6540 : data = 8'h00;
 6541 : data = 8'h00;
 6542 : data = 8'h00;
 6543 : data = 8'h00;
 6544 : data = 8'h00;
 6545 : data = 8'h00;
 6546 : data = 8'h00;
 6547 : data = 8'h00;
 6548 : data = 8'h00;
 6549 : data = 8'h00;
 6550 : data = 8'h00;
 6551 : data = 8'h00;
 6552 : data = 8'h00;
 6553 : data = 8'h00;
 6554 : data = 8'h00;
 6555 : data = 8'h00;
 6556 : data = 8'h00;
 6557 : data = 8'h00;
 6558 : data = 8'h00;
 6559 : data = 8'h00;
 6560 : data = 8'h00;
 6561 : data = 8'h00;
 6562 : data = 8'h00;
 6563 : data = 8'h00;
 6564 : data = 8'h00;
 6565 : data = 8'h00;
 6566 : data = 8'h00;
 6567 : data = 8'h00;
 6568 : data = 8'h00;
 6569 : data = 8'h00;
 6570 : data = 8'h00;
 6571 : data = 8'h00;
 6572 : data = 8'h00;
 6573 : data = 8'h00;
 6574 : data = 8'h00;
 6575 : data = 8'h00;
 6576 : data = 8'h00;
 6577 : data = 8'h00;
 6578 : data = 8'h00;
 6579 : data = 8'h00;
 6580 : data = 8'h00;
 6581 : data = 8'h00;
 6582 : data = 8'h00;
 6583 : data = 8'h00;
 6584 : data = 8'h00;
 6585 : data = 8'h00;
 6586 : data = 8'h00;
 6587 : data = 8'h00;
 6588 : data = 8'h00;
 6589 : data = 8'h00;
 6590 : data = 8'h00;
 6591 : data = 8'h00;
 6592 : data = 8'h00;
 6593 : data = 8'h00;
 6594 : data = 8'h00;
 6595 : data = 8'h00;
 6596 : data = 8'h00;
 6597 : data = 8'h00;
 6598 : data = 8'h00;
 6599 : data = 8'h00;
 6600 : data = 8'h00;
 6601 : data = 8'h00;
 6602 : data = 8'h00;
 6603 : data = 8'h00;
 6604 : data = 8'h00;
 6605 : data = 8'h00;
 6606 : data = 8'h00;
 6607 : data = 8'h00;
 6608 : data = 8'h00;
 6609 : data = 8'h00;
 6610 : data = 8'h00;
 6611 : data = 8'h00;
 6612 : data = 8'h00;
 6613 : data = 8'h00;
 6614 : data = 8'h00;
 6615 : data = 8'h00;
 6616 : data = 8'h00;
 6617 : data = 8'h00;
 6618 : data = 8'h00;
 6619 : data = 8'h00;
 6620 : data = 8'h00;
 6621 : data = 8'h00;
 6622 : data = 8'h00;
 6623 : data = 8'h00;
 6624 : data = 8'h00;
 6625 : data = 8'h00;
 6626 : data = 8'h00;
 6627 : data = 8'h00;
 6628 : data = 8'h00;
 6629 : data = 8'h00;
 6630 : data = 8'h00;
 6631 : data = 8'h00;
 6632 : data = 8'h00;
 6633 : data = 8'h00;
 6634 : data = 8'h00;
 6635 : data = 8'h00;
 6636 : data = 8'h00;
 6637 : data = 8'h00;
 6638 : data = 8'h00;
 6639 : data = 8'h00;
 6640 : data = 8'h00;
 6641 : data = 8'h00;
 6642 : data = 8'h00;
 6643 : data = 8'h00;
 6644 : data = 8'h00;
 6645 : data = 8'h00;
 6646 : data = 8'h00;
 6647 : data = 8'h00;
 6648 : data = 8'h00;
 6649 : data = 8'h00;
 6650 : data = 8'h00;
 6651 : data = 8'h00;
 6652 : data = 8'h00;
 6653 : data = 8'h00;
 6654 : data = 8'h00;
 6655 : data = 8'h00;
 6656 : data = 8'h00;
 6657 : data = 8'h00;
 6658 : data = 8'h00;
 6659 : data = 8'h00;
 6660 : data = 8'h00;
 6661 : data = 8'h00;
 6662 : data = 8'h00;
 6663 : data = 8'h00;
 6664 : data = 8'h00;
 6665 : data = 8'h00;
 6666 : data = 8'h00;
 6667 : data = 8'h00;
 6668 : data = 8'h00;
 6669 : data = 8'h00;
 6670 : data = 8'h00;
 6671 : data = 8'h00;
 6672 : data = 8'h00;
 6673 : data = 8'h00;
 6674 : data = 8'h00;
 6675 : data = 8'h00;
 6676 : data = 8'h00;
 6677 : data = 8'h00;
 6678 : data = 8'h00;
 6679 : data = 8'h00;
 6680 : data = 8'h00;
 6681 : data = 8'h00;
 6682 : data = 8'h00;
 6683 : data = 8'h00;
 6684 : data = 8'h00;
 6685 : data = 8'h00;
 6686 : data = 8'h00;
 6687 : data = 8'h00;
 6688 : data = 8'h00;
 6689 : data = 8'h00;
 6690 : data = 8'h00;
 6691 : data = 8'h00;
 6692 : data = 8'h00;
 6693 : data = 8'h00;
 6694 : data = 8'h00;
 6695 : data = 8'h00;
 6696 : data = 8'h00;
 6697 : data = 8'h00;
 6698 : data = 8'h00;
 6699 : data = 8'h00;
 6700 : data = 8'h00;
 6701 : data = 8'h00;
 6702 : data = 8'h00;
 6703 : data = 8'h00;
 6704 : data = 8'h00;
 6705 : data = 8'h00;
 6706 : data = 8'h00;
 6707 : data = 8'h00;
 6708 : data = 8'h00;
 6709 : data = 8'h00;
 6710 : data = 8'h00;
 6711 : data = 8'h00;
 6712 : data = 8'h00;
 6713 : data = 8'h00;
 6714 : data = 8'h00;
 6715 : data = 8'h00;
 6716 : data = 8'h00;
 6717 : data = 8'h00;
 6718 : data = 8'h00;
 6719 : data = 8'h00;
 6720 : data = 8'h00;
 6721 : data = 8'h00;
 6722 : data = 8'h00;
 6723 : data = 8'h00;
 6724 : data = 8'h00;
 6725 : data = 8'h00;
 6726 : data = 8'h00;
 6727 : data = 8'h00;
 6728 : data = 8'h00;
 6729 : data = 8'h00;
 6730 : data = 8'h00;
 6731 : data = 8'h00;
 6732 : data = 8'h00;
 6733 : data = 8'h00;
 6734 : data = 8'h00;
 6735 : data = 8'h00;
 6736 : data = 8'h00;
 6737 : data = 8'h00;
 6738 : data = 8'h00;
 6739 : data = 8'h00;
 6740 : data = 8'h00;
 6741 : data = 8'h00;
 6742 : data = 8'h00;
 6743 : data = 8'h00;
 6744 : data = 8'h00;
 6745 : data = 8'h00;
 6746 : data = 8'h00;
 6747 : data = 8'h00;
 6748 : data = 8'h00;
 6749 : data = 8'h00;
 6750 : data = 8'h00;
 6751 : data = 8'h00;
 6752 : data = 8'h00;
 6753 : data = 8'h00;
 6754 : data = 8'h00;
 6755 : data = 8'h00;
 6756 : data = 8'h00;
 6757 : data = 8'h00;
 6758 : data = 8'h00;
 6759 : data = 8'h00;
 6760 : data = 8'h00;
 6761 : data = 8'h00;
 6762 : data = 8'h00;
 6763 : data = 8'h00;
 6764 : data = 8'h00;
 6765 : data = 8'h00;
 6766 : data = 8'h00;
 6767 : data = 8'h00;
 6768 : data = 8'h00;
 6769 : data = 8'h00;
 6770 : data = 8'h00;
 6771 : data = 8'h00;
 6772 : data = 8'h00;
 6773 : data = 8'h00;
 6774 : data = 8'h00;
 6775 : data = 8'h00;
 6776 : data = 8'h00;
 6777 : data = 8'h00;
 6778 : data = 8'h00;
 6779 : data = 8'h00;
 6780 : data = 8'h00;
 6781 : data = 8'h00;
 6782 : data = 8'h00;
 6783 : data = 8'h00;
 6784 : data = 8'h00;
 6785 : data = 8'h00;
 6786 : data = 8'h00;
 6787 : data = 8'h00;
 6788 : data = 8'h00;
 6789 : data = 8'h00;
 6790 : data = 8'h00;
 6791 : data = 8'h00;
 6792 : data = 8'h00;
 6793 : data = 8'h00;
 6794 : data = 8'h00;
 6795 : data = 8'h00;
 6796 : data = 8'h00;
 6797 : data = 8'h00;
 6798 : data = 8'h00;
 6799 : data = 8'h00;
 6800 : data = 8'h00;
 6801 : data = 8'h00;
 6802 : data = 8'h00;
 6803 : data = 8'h00;
 6804 : data = 8'h00;
 6805 : data = 8'h00;
 6806 : data = 8'h00;
 6807 : data = 8'h00;
 6808 : data = 8'h00;
 6809 : data = 8'h00;
 6810 : data = 8'h00;
 6811 : data = 8'h00;
 6812 : data = 8'h00;
 6813 : data = 8'h00;
 6814 : data = 8'h00;
 6815 : data = 8'h00;
 6816 : data = 8'h00;
 6817 : data = 8'h00;
 6818 : data = 8'h00;
 6819 : data = 8'h00;
 6820 : data = 8'h00;
 6821 : data = 8'h00;
 6822 : data = 8'h00;
 6823 : data = 8'h00;
 6824 : data = 8'h00;
 6825 : data = 8'h00;
 6826 : data = 8'h00;
 6827 : data = 8'h00;
 6828 : data = 8'h00;
 6829 : data = 8'h00;
 6830 : data = 8'h00;
 6831 : data = 8'h00;
 6832 : data = 8'h00;
 6833 : data = 8'h00;
 6834 : data = 8'h00;
 6835 : data = 8'h00;
 6836 : data = 8'h00;
 6837 : data = 8'h00;
 6838 : data = 8'h00;
 6839 : data = 8'h00;
 6840 : data = 8'h00;
 6841 : data = 8'h00;
 6842 : data = 8'h00;
 6843 : data = 8'h00;
 6844 : data = 8'h00;
 6845 : data = 8'h00;
 6846 : data = 8'h00;
 6847 : data = 8'h00;
 6848 : data = 8'h00;
 6849 : data = 8'h00;
 6850 : data = 8'h00;
 6851 : data = 8'h00;
 6852 : data = 8'h00;
 6853 : data = 8'h00;
 6854 : data = 8'h00;
 6855 : data = 8'h00;
 6856 : data = 8'h00;
 6857 : data = 8'h00;
 6858 : data = 8'h00;
 6859 : data = 8'h00;
 6860 : data = 8'h00;
 6861 : data = 8'h00;
 6862 : data = 8'h00;
 6863 : data = 8'h00;
 6864 : data = 8'h00;
 6865 : data = 8'h00;
 6866 : data = 8'h00;
 6867 : data = 8'h00;
 6868 : data = 8'h00;
 6869 : data = 8'h00;
 6870 : data = 8'h00;
 6871 : data = 8'h00;
 6872 : data = 8'h00;
 6873 : data = 8'h00;
 6874 : data = 8'h00;
 6875 : data = 8'h00;
 6876 : data = 8'h00;
 6877 : data = 8'h00;
 6878 : data = 8'h00;
 6879 : data = 8'h00;
 6880 : data = 8'h00;
 6881 : data = 8'h00;
 6882 : data = 8'h00;
 6883 : data = 8'h00;
 6884 : data = 8'h00;
 6885 : data = 8'h00;
 6886 : data = 8'h00;
 6887 : data = 8'h00;
 6888 : data = 8'h00;
 6889 : data = 8'h00;
 6890 : data = 8'h00;
 6891 : data = 8'h00;
 6892 : data = 8'h00;
 6893 : data = 8'h00;
 6894 : data = 8'h00;
 6895 : data = 8'h00;
 6896 : data = 8'h00;
 6897 : data = 8'h00;
 6898 : data = 8'h00;
 6899 : data = 8'h00;
 6900 : data = 8'h00;
 6901 : data = 8'h00;
 6902 : data = 8'h00;
 6903 : data = 8'h00;
 6904 : data = 8'h00;
 6905 : data = 8'h00;
 6906 : data = 8'h00;
 6907 : data = 8'h00;
 6908 : data = 8'h00;
 6909 : data = 8'h00;
 6910 : data = 8'h00;
 6911 : data = 8'h00;
 6912 : data = 8'h00;
 6913 : data = 8'h00;
 6914 : data = 8'h00;
 6915 : data = 8'h00;
 6916 : data = 8'h00;
 6917 : data = 8'h00;
 6918 : data = 8'h00;
 6919 : data = 8'h00;
 6920 : data = 8'h00;
 6921 : data = 8'h00;
 6922 : data = 8'h00;
 6923 : data = 8'h00;
 6924 : data = 8'h00;
 6925 : data = 8'h00;
 6926 : data = 8'h00;
 6927 : data = 8'h00;
 6928 : data = 8'h00;
 6929 : data = 8'h00;
 6930 : data = 8'h00;
 6931 : data = 8'h00;
 6932 : data = 8'h00;
 6933 : data = 8'h00;
 6934 : data = 8'h00;
 6935 : data = 8'h00;
 6936 : data = 8'h00;
 6937 : data = 8'h00;
 6938 : data = 8'h00;
 6939 : data = 8'h00;
 6940 : data = 8'h00;
 6941 : data = 8'h00;
 6942 : data = 8'h00;
 6943 : data = 8'h00;
 6944 : data = 8'h00;
 6945 : data = 8'h00;
 6946 : data = 8'h00;
 6947 : data = 8'h00;
 6948 : data = 8'h00;
 6949 : data = 8'h00;
 6950 : data = 8'h00;
 6951 : data = 8'h00;
 6952 : data = 8'h00;
 6953 : data = 8'h00;
 6954 : data = 8'h00;
 6955 : data = 8'h00;
 6956 : data = 8'h00;
 6957 : data = 8'h00;
 6958 : data = 8'h00;
 6959 : data = 8'h00;
 6960 : data = 8'h00;
 6961 : data = 8'h00;
 6962 : data = 8'h00;
 6963 : data = 8'h00;
 6964 : data = 8'h00;
 6965 : data = 8'h00;
 6966 : data = 8'h00;
 6967 : data = 8'h00;
 6968 : data = 8'h00;
 6969 : data = 8'h00;
 6970 : data = 8'h00;
 6971 : data = 8'h00;
 6972 : data = 8'h00;
 6973 : data = 8'h00;
 6974 : data = 8'h00;
 6975 : data = 8'h00;
 6976 : data = 8'h00;
 6977 : data = 8'h00;
 6978 : data = 8'h00;
 6979 : data = 8'h00;
 6980 : data = 8'h00;
 6981 : data = 8'h00;
 6982 : data = 8'h00;
 6983 : data = 8'h00;
 6984 : data = 8'h00;
 6985 : data = 8'h00;
 6986 : data = 8'h00;
 6987 : data = 8'h00;
 6988 : data = 8'h00;
 6989 : data = 8'h00;
 6990 : data = 8'h00;
 6991 : data = 8'h00;
 6992 : data = 8'h00;
 6993 : data = 8'h00;
 6994 : data = 8'h00;
 6995 : data = 8'h00;
 6996 : data = 8'h00;
 6997 : data = 8'h00;
 6998 : data = 8'h00;
 6999 : data = 8'h00;
 7000 : data = 8'h00;
 7001 : data = 8'h00;
 7002 : data = 8'h00;
 7003 : data = 8'h00;
 7004 : data = 8'h00;
 7005 : data = 8'h00;
 7006 : data = 8'h00;
 7007 : data = 8'h00;
 7008 : data = 8'h00;
 7009 : data = 8'h00;
 7010 : data = 8'h00;
 7011 : data = 8'h00;
 7012 : data = 8'h00;
 7013 : data = 8'h00;
 7014 : data = 8'h00;
 7015 : data = 8'h00;
 7016 : data = 8'h00;
 7017 : data = 8'h00;
 7018 : data = 8'h00;
 7019 : data = 8'h00;
 7020 : data = 8'h00;
 7021 : data = 8'h00;
 7022 : data = 8'h00;
 7023 : data = 8'h00;
 7024 : data = 8'h00;
 7025 : data = 8'h00;
 7026 : data = 8'h00;
 7027 : data = 8'h00;
 7028 : data = 8'h00;
 7029 : data = 8'h00;
 7030 : data = 8'h00;
 7031 : data = 8'h00;
 7032 : data = 8'h00;
 7033 : data = 8'h00;
 7034 : data = 8'h00;
 7035 : data = 8'h00;
 7036 : data = 8'h00;
 7037 : data = 8'h00;
 7038 : data = 8'h00;
 7039 : data = 8'h00;
 7040 : data = 8'h00;
 7041 : data = 8'h00;
 7042 : data = 8'h00;
 7043 : data = 8'h00;
 7044 : data = 8'h00;
 7045 : data = 8'h00;
 7046 : data = 8'h00;
 7047 : data = 8'h00;
 7048 : data = 8'h00;
 7049 : data = 8'h00;
 7050 : data = 8'h00;
 7051 : data = 8'h00;
 7052 : data = 8'h00;
 7053 : data = 8'h00;
 7054 : data = 8'h00;
 7055 : data = 8'h00;
 7056 : data = 8'h00;
 7057 : data = 8'h00;
 7058 : data = 8'h00;
 7059 : data = 8'h00;
 7060 : data = 8'h00;
 7061 : data = 8'h00;
 7062 : data = 8'h00;
 7063 : data = 8'h00;
 7064 : data = 8'h00;
 7065 : data = 8'h00;
 7066 : data = 8'h00;
 7067 : data = 8'h00;
 7068 : data = 8'h00;
 7069 : data = 8'h00;
 7070 : data = 8'h00;
 7071 : data = 8'h00;
 7072 : data = 8'h00;
 7073 : data = 8'h00;
 7074 : data = 8'h00;
 7075 : data = 8'h00;
 7076 : data = 8'h00;
 7077 : data = 8'h00;
 7078 : data = 8'h00;
 7079 : data = 8'h00;
 7080 : data = 8'h00;
 7081 : data = 8'h00;
 7082 : data = 8'h00;
 7083 : data = 8'h00;
 7084 : data = 8'h00;
 7085 : data = 8'h00;
 7086 : data = 8'h00;
 7087 : data = 8'h00;
 7088 : data = 8'h00;
 7089 : data = 8'h00;
 7090 : data = 8'h00;
 7091 : data = 8'h00;
 7092 : data = 8'h00;
 7093 : data = 8'h00;
 7094 : data = 8'h00;
 7095 : data = 8'h00;
 7096 : data = 8'h00;
 7097 : data = 8'h00;
 7098 : data = 8'h00;
 7099 : data = 8'h00;
 7100 : data = 8'h00;
 7101 : data = 8'h00;
 7102 : data = 8'h00;
 7103 : data = 8'h00;
 7104 : data = 8'h00;
 7105 : data = 8'h00;
 7106 : data = 8'h00;
 7107 : data = 8'h00;
 7108 : data = 8'h00;
 7109 : data = 8'h00;
 7110 : data = 8'h00;
 7111 : data = 8'h00;
 7112 : data = 8'h00;
 7113 : data = 8'h00;
 7114 : data = 8'h00;
 7115 : data = 8'h00;
 7116 : data = 8'h00;
 7117 : data = 8'h00;
 7118 : data = 8'h00;
 7119 : data = 8'h00;
 7120 : data = 8'h00;
 7121 : data = 8'h00;
 7122 : data = 8'h00;
 7123 : data = 8'h00;
 7124 : data = 8'h00;
 7125 : data = 8'h00;
 7126 : data = 8'h00;
 7127 : data = 8'h00;
 7128 : data = 8'h00;
 7129 : data = 8'h00;
 7130 : data = 8'h00;
 7131 : data = 8'h00;
 7132 : data = 8'h00;
 7133 : data = 8'h00;
 7134 : data = 8'h00;
 7135 : data = 8'h00;
 7136 : data = 8'h00;
 7137 : data = 8'h00;
 7138 : data = 8'h00;
 7139 : data = 8'h00;
 7140 : data = 8'h00;
 7141 : data = 8'h00;
 7142 : data = 8'h00;
 7143 : data = 8'h00;
 7144 : data = 8'h00;
 7145 : data = 8'h00;
 7146 : data = 8'h00;
 7147 : data = 8'h00;
 7148 : data = 8'h00;
 7149 : data = 8'h00;
 7150 : data = 8'h00;
 7151 : data = 8'h00;
 7152 : data = 8'h00;
 7153 : data = 8'h00;
 7154 : data = 8'h00;
 7155 : data = 8'h00;
 7156 : data = 8'h00;
 7157 : data = 8'h00;
 7158 : data = 8'h00;
 7159 : data = 8'h00;
 7160 : data = 8'h00;
 7161 : data = 8'h00;
 7162 : data = 8'h00;
 7163 : data = 8'h00;
 7164 : data = 8'h00;
 7165 : data = 8'h00;
 7166 : data = 8'h00;
 7167 : data = 8'h00;
 7168 : data = 8'h00;
 7169 : data = 8'h00;
 7170 : data = 8'h00;
 7171 : data = 8'h00;
 7172 : data = 8'h00;
 7173 : data = 8'h00;
 7174 : data = 8'h00;
 7175 : data = 8'h00;
 7176 : data = 8'h00;
 7177 : data = 8'h00;
 7178 : data = 8'h00;
 7179 : data = 8'h00;
 7180 : data = 8'h00;
 7181 : data = 8'h00;
 7182 : data = 8'h00;
 7183 : data = 8'h00;
 7184 : data = 8'h00;
 7185 : data = 8'h00;
 7186 : data = 8'h00;
 7187 : data = 8'h00;
 7188 : data = 8'h00;
 7189 : data = 8'h00;
 7190 : data = 8'h00;
 7191 : data = 8'h00;
 7192 : data = 8'h00;
 7193 : data = 8'h00;
 7194 : data = 8'h00;
 7195 : data = 8'h00;
 7196 : data = 8'h00;
 7197 : data = 8'h00;
 7198 : data = 8'h00;
 7199 : data = 8'h00;
 7200 : data = 8'h00;
 7201 : data = 8'h00;
 7202 : data = 8'h00;
 7203 : data = 8'h00;
 7204 : data = 8'h00;
 7205 : data = 8'h00;
 7206 : data = 8'h00;
 7207 : data = 8'h00;
 7208 : data = 8'h00;
 7209 : data = 8'h00;
 7210 : data = 8'h00;
 7211 : data = 8'h00;
 7212 : data = 8'h00;
 7213 : data = 8'h00;
 7214 : data = 8'h00;
 7215 : data = 8'h00;
 7216 : data = 8'h00;
 7217 : data = 8'h00;
 7218 : data = 8'h00;
 7219 : data = 8'h00;
 7220 : data = 8'h00;
 7221 : data = 8'h00;
 7222 : data = 8'h00;
 7223 : data = 8'h00;
 7224 : data = 8'h00;
 7225 : data = 8'h00;
 7226 : data = 8'h00;
 7227 : data = 8'h00;
 7228 : data = 8'h00;
 7229 : data = 8'h00;
 7230 : data = 8'h00;
 7231 : data = 8'h00;
 7232 : data = 8'h00;
 7233 : data = 8'h00;
 7234 : data = 8'h00;
 7235 : data = 8'h00;
 7236 : data = 8'h00;
 7237 : data = 8'h00;
 7238 : data = 8'h00;
 7239 : data = 8'h00;
 7240 : data = 8'h00;
 7241 : data = 8'h00;
 7242 : data = 8'h00;
 7243 : data = 8'h00;
 7244 : data = 8'h00;
 7245 : data = 8'h00;
 7246 : data = 8'h00;
 7247 : data = 8'h00;
 7248 : data = 8'h00;
 7249 : data = 8'h00;
 7250 : data = 8'h00;
 7251 : data = 8'h00;
 7252 : data = 8'h00;
 7253 : data = 8'h00;
 7254 : data = 8'h00;
 7255 : data = 8'h00;
 7256 : data = 8'h00;
 7257 : data = 8'h00;
 7258 : data = 8'h00;
 7259 : data = 8'h00;
 7260 : data = 8'h00;
 7261 : data = 8'h00;
 7262 : data = 8'h00;
 7263 : data = 8'h00;
 7264 : data = 8'h00;
 7265 : data = 8'h00;
 7266 : data = 8'h00;
 7267 : data = 8'h00;
 7268 : data = 8'h00;
 7269 : data = 8'h00;
 7270 : data = 8'h00;
 7271 : data = 8'h00;
 7272 : data = 8'h00;
 7273 : data = 8'h00;
 7274 : data = 8'h00;
 7275 : data = 8'h00;
 7276 : data = 8'h00;
 7277 : data = 8'h00;
 7278 : data = 8'h00;
 7279 : data = 8'h00;
 7280 : data = 8'h00;
 7281 : data = 8'h00;
 7282 : data = 8'h00;
 7283 : data = 8'h00;
 7284 : data = 8'h00;
 7285 : data = 8'h00;
 7286 : data = 8'h00;
 7287 : data = 8'h00;
 7288 : data = 8'h00;
 7289 : data = 8'h00;
 7290 : data = 8'h00;
 7291 : data = 8'h00;
 7292 : data = 8'h00;
 7293 : data = 8'h00;
 7294 : data = 8'h00;
 7295 : data = 8'h00;
 7296 : data = 8'h00;
 7297 : data = 8'h00;
 7298 : data = 8'h00;
 7299 : data = 8'h00;
 7300 : data = 8'h00;
 7301 : data = 8'h00;
 7302 : data = 8'h00;
 7303 : data = 8'h00;
 7304 : data = 8'h00;
 7305 : data = 8'h00;
 7306 : data = 8'h00;
 7307 : data = 8'h00;
 7308 : data = 8'h00;
 7309 : data = 8'h00;
 7310 : data = 8'h00;
 7311 : data = 8'h00;
 7312 : data = 8'h00;
 7313 : data = 8'h00;
 7314 : data = 8'h00;
 7315 : data = 8'h00;
 7316 : data = 8'h00;
 7317 : data = 8'h00;
 7318 : data = 8'h00;
 7319 : data = 8'h00;
 7320 : data = 8'h00;
 7321 : data = 8'h00;
 7322 : data = 8'h00;
 7323 : data = 8'h00;
 7324 : data = 8'h00;
 7325 : data = 8'h00;
 7326 : data = 8'h00;
 7327 : data = 8'h00;
 7328 : data = 8'h00;
 7329 : data = 8'h00;
 7330 : data = 8'h00;
 7331 : data = 8'h00;
 7332 : data = 8'h00;
 7333 : data = 8'h00;
 7334 : data = 8'h00;
 7335 : data = 8'h00;
 7336 : data = 8'h00;
 7337 : data = 8'h00;
 7338 : data = 8'h00;
 7339 : data = 8'h00;
 7340 : data = 8'h00;
 7341 : data = 8'h00;
 7342 : data = 8'h00;
 7343 : data = 8'h00;
 7344 : data = 8'h00;
 7345 : data = 8'h00;
 7346 : data = 8'h00;
 7347 : data = 8'h00;
 7348 : data = 8'h00;
 7349 : data = 8'h00;
 7350 : data = 8'h00;
 7351 : data = 8'h00;
 7352 : data = 8'h00;
 7353 : data = 8'h00;
 7354 : data = 8'h00;
 7355 : data = 8'h00;
 7356 : data = 8'h00;
 7357 : data = 8'h00;
 7358 : data = 8'h00;
 7359 : data = 8'h00;
 7360 : data = 8'h00;
 7361 : data = 8'h00;
 7362 : data = 8'h00;
 7363 : data = 8'h00;
 7364 : data = 8'h00;
 7365 : data = 8'h00;
 7366 : data = 8'h00;
 7367 : data = 8'h00;
 7368 : data = 8'h00;
 7369 : data = 8'h00;
 7370 : data = 8'h00;
 7371 : data = 8'h00;
 7372 : data = 8'h00;
 7373 : data = 8'h00;
 7374 : data = 8'h00;
 7375 : data = 8'h00;
 7376 : data = 8'h00;
 7377 : data = 8'h00;
 7378 : data = 8'h00;
 7379 : data = 8'h00;
 7380 : data = 8'h00;
 7381 : data = 8'h00;
 7382 : data = 8'h00;
 7383 : data = 8'h00;
 7384 : data = 8'h00;
 7385 : data = 8'h00;
 7386 : data = 8'h00;
 7387 : data = 8'h00;
 7388 : data = 8'h00;
 7389 : data = 8'h00;
 7390 : data = 8'h00;
 7391 : data = 8'h00;
 7392 : data = 8'h00;
 7393 : data = 8'h00;
 7394 : data = 8'h00;
 7395 : data = 8'h00;
 7396 : data = 8'h00;
 7397 : data = 8'h00;
 7398 : data = 8'h00;
 7399 : data = 8'h00;
 7400 : data = 8'h00;
 7401 : data = 8'h00;
 7402 : data = 8'h00;
 7403 : data = 8'h00;
 7404 : data = 8'h00;
 7405 : data = 8'h00;
 7406 : data = 8'h00;
 7407 : data = 8'h00;
 7408 : data = 8'h00;
 7409 : data = 8'h00;
 7410 : data = 8'h00;
 7411 : data = 8'h00;
 7412 : data = 8'h00;
 7413 : data = 8'h00;
 7414 : data = 8'h00;
 7415 : data = 8'h00;
 7416 : data = 8'h00;
 7417 : data = 8'h00;
 7418 : data = 8'h00;
 7419 : data = 8'h00;
 7420 : data = 8'h00;
 7421 : data = 8'h00;
 7422 : data = 8'h00;
 7423 : data = 8'h00;
 7424 : data = 8'h00;
 7425 : data = 8'h00;
 7426 : data = 8'h00;
 7427 : data = 8'h00;
 7428 : data = 8'h00;
 7429 : data = 8'h00;
 7430 : data = 8'h00;
 7431 : data = 8'h00;
 7432 : data = 8'h00;
 7433 : data = 8'h00;
 7434 : data = 8'h00;
 7435 : data = 8'h00;
 7436 : data = 8'h00;
 7437 : data = 8'h00;
 7438 : data = 8'h00;
 7439 : data = 8'h00;
 7440 : data = 8'h00;
 7441 : data = 8'h00;
 7442 : data = 8'h00;
 7443 : data = 8'h00;
 7444 : data = 8'h00;
 7445 : data = 8'h00;
 7446 : data = 8'h00;
 7447 : data = 8'h00;
 7448 : data = 8'h00;
 7449 : data = 8'h00;
 7450 : data = 8'h00;
 7451 : data = 8'h00;
 7452 : data = 8'h00;
 7453 : data = 8'h00;
 7454 : data = 8'h00;
 7455 : data = 8'h00;
 7456 : data = 8'h00;
 7457 : data = 8'h00;
 7458 : data = 8'h00;
 7459 : data = 8'h00;
 7460 : data = 8'h00;
 7461 : data = 8'h00;
 7462 : data = 8'h00;
 7463 : data = 8'h00;
 7464 : data = 8'h00;
 7465 : data = 8'h00;
 7466 : data = 8'h00;
 7467 : data = 8'h00;
 7468 : data = 8'h00;
 7469 : data = 8'h00;
 7470 : data = 8'h00;
 7471 : data = 8'h00;
 7472 : data = 8'h00;
 7473 : data = 8'h00;
 7474 : data = 8'h00;
 7475 : data = 8'h00;
 7476 : data = 8'h00;
 7477 : data = 8'h00;
 7478 : data = 8'h00;
 7479 : data = 8'h00;
 7480 : data = 8'h00;
 7481 : data = 8'h00;
 7482 : data = 8'h00;
 7483 : data = 8'h00;
 7484 : data = 8'h00;
 7485 : data = 8'h00;
 7486 : data = 8'h00;
 7487 : data = 8'h00;
 7488 : data = 8'h00;
 7489 : data = 8'h00;
 7490 : data = 8'h00;
 7491 : data = 8'h00;
 7492 : data = 8'h00;
 7493 : data = 8'h00;
 7494 : data = 8'h00;
 7495 : data = 8'h00;
 7496 : data = 8'h00;
 7497 : data = 8'h00;
 7498 : data = 8'h00;
 7499 : data = 8'h00;
 7500 : data = 8'h00;
 7501 : data = 8'h00;
 7502 : data = 8'h00;
 7503 : data = 8'h00;
 7504 : data = 8'h00;
 7505 : data = 8'h00;
 7506 : data = 8'h00;
 7507 : data = 8'h00;
 7508 : data = 8'h00;
 7509 : data = 8'h00;
 7510 : data = 8'h00;
 7511 : data = 8'h00;
 7512 : data = 8'h00;
 7513 : data = 8'h00;
 7514 : data = 8'h00;
 7515 : data = 8'h00;
 7516 : data = 8'h00;
 7517 : data = 8'h00;
 7518 : data = 8'h00;
 7519 : data = 8'h00;
 7520 : data = 8'h00;
 7521 : data = 8'h00;
 7522 : data = 8'h00;
 7523 : data = 8'h00;
 7524 : data = 8'h00;
 7525 : data = 8'h00;
 7526 : data = 8'h00;
 7527 : data = 8'h00;
 7528 : data = 8'h00;
 7529 : data = 8'h00;
 7530 : data = 8'h00;
 7531 : data = 8'h00;
 7532 : data = 8'h00;
 7533 : data = 8'h00;
 7534 : data = 8'h00;
 7535 : data = 8'h00;
 7536 : data = 8'h00;
 7537 : data = 8'h00;
 7538 : data = 8'h00;
 7539 : data = 8'h00;
 7540 : data = 8'h00;
 7541 : data = 8'h00;
 7542 : data = 8'h00;
 7543 : data = 8'h00;
 7544 : data = 8'h00;
 7545 : data = 8'h00;
 7546 : data = 8'h00;
 7547 : data = 8'h00;
 7548 : data = 8'h00;
 7549 : data = 8'h00;
 7550 : data = 8'h00;
 7551 : data = 8'h00;
 7552 : data = 8'h00;
 7553 : data = 8'h00;
 7554 : data = 8'h00;
 7555 : data = 8'h00;
 7556 : data = 8'h00;
 7557 : data = 8'h00;
 7558 : data = 8'h00;
 7559 : data = 8'h00;
 7560 : data = 8'h00;
 7561 : data = 8'h00;
 7562 : data = 8'h00;
 7563 : data = 8'h00;
 7564 : data = 8'h00;
 7565 : data = 8'h00;
 7566 : data = 8'h00;
 7567 : data = 8'h00;
 7568 : data = 8'h00;
 7569 : data = 8'h00;
 7570 : data = 8'h00;
 7571 : data = 8'h00;
 7572 : data = 8'h00;
 7573 : data = 8'h00;
 7574 : data = 8'h00;
 7575 : data = 8'h00;
 7576 : data = 8'h00;
 7577 : data = 8'h00;
 7578 : data = 8'h00;
 7579 : data = 8'h00;
 7580 : data = 8'h00;
 7581 : data = 8'h00;
 7582 : data = 8'h00;
 7583 : data = 8'h00;
 7584 : data = 8'h00;
 7585 : data = 8'h00;
 7586 : data = 8'h00;
 7587 : data = 8'h00;
 7588 : data = 8'h00;
 7589 : data = 8'h00;
 7590 : data = 8'h00;
 7591 : data = 8'h00;
 7592 : data = 8'h00;
 7593 : data = 8'h00;
 7594 : data = 8'h00;
 7595 : data = 8'h00;
 7596 : data = 8'h00;
 7597 : data = 8'h00;
 7598 : data = 8'h00;
 7599 : data = 8'h00;
 7600 : data = 8'h00;
 7601 : data = 8'h00;
 7602 : data = 8'h00;
 7603 : data = 8'h00;
 7604 : data = 8'h00;
 7605 : data = 8'h00;
 7606 : data = 8'h00;
 7607 : data = 8'h00;
 7608 : data = 8'h00;
 7609 : data = 8'h00;
 7610 : data = 8'h00;
 7611 : data = 8'h00;
 7612 : data = 8'h00;
 7613 : data = 8'h00;
 7614 : data = 8'h00;
 7615 : data = 8'h00;
 7616 : data = 8'h00;
 7617 : data = 8'h00;
 7618 : data = 8'h00;
 7619 : data = 8'h00;
 7620 : data = 8'h00;
 7621 : data = 8'h00;
 7622 : data = 8'h00;
 7623 : data = 8'h00;
 7624 : data = 8'h00;
 7625 : data = 8'h00;
 7626 : data = 8'h00;
 7627 : data = 8'h00;
 7628 : data = 8'h00;
 7629 : data = 8'h00;
 7630 : data = 8'h00;
 7631 : data = 8'h00;
 7632 : data = 8'h00;
 7633 : data = 8'h00;
 7634 : data = 8'h00;
 7635 : data = 8'h00;
 7636 : data = 8'h00;
 7637 : data = 8'h00;
 7638 : data = 8'h00;
 7639 : data = 8'h00;
 7640 : data = 8'h00;
 7641 : data = 8'h00;
 7642 : data = 8'h00;
 7643 : data = 8'h00;
 7644 : data = 8'h00;
 7645 : data = 8'h00;
 7646 : data = 8'h00;
 7647 : data = 8'h00;
 7648 : data = 8'h00;
 7649 : data = 8'h00;
 7650 : data = 8'h00;
 7651 : data = 8'h00;
 7652 : data = 8'h00;
 7653 : data = 8'h00;
 7654 : data = 8'h00;
 7655 : data = 8'h00;
 7656 : data = 8'h00;
 7657 : data = 8'h00;
 7658 : data = 8'h00;
 7659 : data = 8'h00;
 7660 : data = 8'h00;
 7661 : data = 8'h00;
 7662 : data = 8'h00;
 7663 : data = 8'h00;
 7664 : data = 8'h00;
 7665 : data = 8'h00;
 7666 : data = 8'h00;
 7667 : data = 8'h00;
 7668 : data = 8'h00;
 7669 : data = 8'h00;
 7670 : data = 8'h00;
 7671 : data = 8'h00;
 7672 : data = 8'h00;
 7673 : data = 8'h00;
 7674 : data = 8'h00;
 7675 : data = 8'h00;
 7676 : data = 8'h00;
 7677 : data = 8'h00;
 7678 : data = 8'h00;
 7679 : data = 8'h00;
 7680 : data = 8'h00;
 7681 : data = 8'h00;
 7682 : data = 8'h00;
 7683 : data = 8'h00;
 7684 : data = 8'h00;
 7685 : data = 8'h00;
 7686 : data = 8'h00;
 7687 : data = 8'h00;
 7688 : data = 8'h00;
 7689 : data = 8'h00;
 7690 : data = 8'h00;
 7691 : data = 8'h00;
 7692 : data = 8'h00;
 7693 : data = 8'h00;
 7694 : data = 8'h00;
 7695 : data = 8'h00;
 7696 : data = 8'h00;
 7697 : data = 8'h00;
 7698 : data = 8'h00;
 7699 : data = 8'h00;
 7700 : data = 8'h00;
 7701 : data = 8'h00;
 7702 : data = 8'h00;
 7703 : data = 8'h00;
 7704 : data = 8'h00;
 7705 : data = 8'h00;
 7706 : data = 8'h00;
 7707 : data = 8'h00;
 7708 : data = 8'h00;
 7709 : data = 8'h00;
 7710 : data = 8'h00;
 7711 : data = 8'h00;
 7712 : data = 8'h00;
 7713 : data = 8'h00;
 7714 : data = 8'h00;
 7715 : data = 8'h00;
 7716 : data = 8'h00;
 7717 : data = 8'h00;
 7718 : data = 8'h00;
 7719 : data = 8'h00;
 7720 : data = 8'h00;
 7721 : data = 8'h00;
 7722 : data = 8'h00;
 7723 : data = 8'h00;
 7724 : data = 8'h00;
 7725 : data = 8'h00;
 7726 : data = 8'h00;
 7727 : data = 8'h00;
 7728 : data = 8'h00;
 7729 : data = 8'h00;
 7730 : data = 8'h00;
 7731 : data = 8'h00;
 7732 : data = 8'h00;
 7733 : data = 8'h00;
 7734 : data = 8'h00;
 7735 : data = 8'h00;
 7736 : data = 8'h00;
 7737 : data = 8'h00;
 7738 : data = 8'h00;
 7739 : data = 8'h00;
 7740 : data = 8'h00;
 7741 : data = 8'h00;
 7742 : data = 8'h00;
 7743 : data = 8'h00;
 7744 : data = 8'h00;
 7745 : data = 8'h00;
 7746 : data = 8'h00;
 7747 : data = 8'h00;
 7748 : data = 8'h00;
 7749 : data = 8'h00;
 7750 : data = 8'h00;
 7751 : data = 8'h00;
 7752 : data = 8'h00;
 7753 : data = 8'h00;
 7754 : data = 8'h00;
 7755 : data = 8'h00;
 7756 : data = 8'h00;
 7757 : data = 8'h00;
 7758 : data = 8'h00;
 7759 : data = 8'h00;
 7760 : data = 8'h00;
 7761 : data = 8'h00;
 7762 : data = 8'h00;
 7763 : data = 8'h00;
 7764 : data = 8'h00;
 7765 : data = 8'h00;
 7766 : data = 8'h00;
 7767 : data = 8'h00;
 7768 : data = 8'h00;
 7769 : data = 8'h00;
 7770 : data = 8'h00;
 7771 : data = 8'h00;
 7772 : data = 8'h00;
 7773 : data = 8'h00;
 7774 : data = 8'h00;
 7775 : data = 8'h00;
 7776 : data = 8'h00;
 7777 : data = 8'h00;
 7778 : data = 8'h00;
 7779 : data = 8'h00;
 7780 : data = 8'h00;
 7781 : data = 8'h00;
 7782 : data = 8'h00;
 7783 : data = 8'h00;
 7784 : data = 8'h00;
 7785 : data = 8'h00;
 7786 : data = 8'h00;
 7787 : data = 8'h00;
 7788 : data = 8'h00;
 7789 : data = 8'h00;
 7790 : data = 8'h00;
 7791 : data = 8'h00;
 7792 : data = 8'h00;
 7793 : data = 8'h00;
 7794 : data = 8'h00;
 7795 : data = 8'h00;
 7796 : data = 8'h00;
 7797 : data = 8'h00;
 7798 : data = 8'h00;
 7799 : data = 8'h00;
 7800 : data = 8'h00;
 7801 : data = 8'h00;
 7802 : data = 8'h00;
 7803 : data = 8'h00;
 7804 : data = 8'h00;
 7805 : data = 8'h00;
 7806 : data = 8'h00;
 7807 : data = 8'h00;
 7808 : data = 8'h00;
 7809 : data = 8'h00;
 7810 : data = 8'h00;
 7811 : data = 8'h00;
 7812 : data = 8'h00;
 7813 : data = 8'h00;
 7814 : data = 8'h00;
 7815 : data = 8'h00;
 7816 : data = 8'h00;
 7817 : data = 8'h00;
 7818 : data = 8'h00;
 7819 : data = 8'h00;
 7820 : data = 8'h00;
 7821 : data = 8'h00;
 7822 : data = 8'h00;
 7823 : data = 8'h00;
 7824 : data = 8'h00;
 7825 : data = 8'h00;
 7826 : data = 8'h00;
 7827 : data = 8'h00;
 7828 : data = 8'h00;
 7829 : data = 8'h00;
 7830 : data = 8'h00;
 7831 : data = 8'h00;
 7832 : data = 8'h00;
 7833 : data = 8'h00;
 7834 : data = 8'h00;
 7835 : data = 8'h00;
 7836 : data = 8'h00;
 7837 : data = 8'h00;
 7838 : data = 8'h00;
 7839 : data = 8'h00;
 7840 : data = 8'h00;
 7841 : data = 8'h00;
 7842 : data = 8'h00;
 7843 : data = 8'h00;
 7844 : data = 8'h00;
 7845 : data = 8'h00;
 7846 : data = 8'h00;
 7847 : data = 8'h00;
 7848 : data = 8'h00;
 7849 : data = 8'h00;
 7850 : data = 8'h00;
 7851 : data = 8'h00;
 7852 : data = 8'h00;
 7853 : data = 8'h00;
 7854 : data = 8'h00;
 7855 : data = 8'h00;
 7856 : data = 8'h00;
 7857 : data = 8'h00;
 7858 : data = 8'h00;
 7859 : data = 8'h00;
 7860 : data = 8'h00;
 7861 : data = 8'h00;
 7862 : data = 8'h00;
 7863 : data = 8'h00;
 7864 : data = 8'h00;
 7865 : data = 8'h00;
 7866 : data = 8'h00;
 7867 : data = 8'h00;
 7868 : data = 8'h00;
 7869 : data = 8'h00;
 7870 : data = 8'h00;
 7871 : data = 8'h00;
 7872 : data = 8'h00;
 7873 : data = 8'h00;
 7874 : data = 8'h00;
 7875 : data = 8'h00;
 7876 : data = 8'h00;
 7877 : data = 8'h00;
 7878 : data = 8'h00;
 7879 : data = 8'h00;
 7880 : data = 8'h00;
 7881 : data = 8'h00;
 7882 : data = 8'h00;
 7883 : data = 8'h00;
 7884 : data = 8'h00;
 7885 : data = 8'h00;
 7886 : data = 8'h00;
 7887 : data = 8'h00;
 7888 : data = 8'h00;
 7889 : data = 8'h00;
 7890 : data = 8'h00;
 7891 : data = 8'h00;
 7892 : data = 8'h00;
 7893 : data = 8'h00;
 7894 : data = 8'h00;
 7895 : data = 8'h00;
 7896 : data = 8'h00;
 7897 : data = 8'h00;
 7898 : data = 8'h00;
 7899 : data = 8'h00;
 7900 : data = 8'h00;
 7901 : data = 8'h00;
 7902 : data = 8'h00;
 7903 : data = 8'h00;
 7904 : data = 8'h00;
 7905 : data = 8'h00;
 7906 : data = 8'h00;
 7907 : data = 8'h00;
 7908 : data = 8'h00;
 7909 : data = 8'h00;
 7910 : data = 8'h00;
 7911 : data = 8'h00;
 7912 : data = 8'h00;
 7913 : data = 8'h00;
 7914 : data = 8'h00;
 7915 : data = 8'h00;
 7916 : data = 8'h00;
 7917 : data = 8'h00;
 7918 : data = 8'h00;
 7919 : data = 8'h00;
 7920 : data = 8'h00;
 7921 : data = 8'h00;
 7922 : data = 8'h00;
 7923 : data = 8'h00;
 7924 : data = 8'h00;
 7925 : data = 8'h00;
 7926 : data = 8'h00;
 7927 : data = 8'h00;
 7928 : data = 8'h00;
 7929 : data = 8'h00;
 7930 : data = 8'h00;
 7931 : data = 8'h00;
 7932 : data = 8'h00;
 7933 : data = 8'h00;
 7934 : data = 8'h00;
 7935 : data = 8'h00;
 7936 : data = 8'h00;
 7937 : data = 8'h00;
 7938 : data = 8'h00;
 7939 : data = 8'h00;
 7940 : data = 8'h00;
 7941 : data = 8'h00;
 7942 : data = 8'h00;
 7943 : data = 8'h00;
 7944 : data = 8'h00;
 7945 : data = 8'h00;
 7946 : data = 8'h00;
 7947 : data = 8'h00;
 7948 : data = 8'h00;
 7949 : data = 8'h00;
 7950 : data = 8'h00;
 7951 : data = 8'h00;
 7952 : data = 8'h00;
 7953 : data = 8'h00;
 7954 : data = 8'h00;
 7955 : data = 8'h00;
 7956 : data = 8'h00;
 7957 : data = 8'h00;
 7958 : data = 8'h00;
 7959 : data = 8'h00;
 7960 : data = 8'h00;
 7961 : data = 8'h00;
 7962 : data = 8'h00;
 7963 : data = 8'h00;
 7964 : data = 8'h00;
 7965 : data = 8'h00;
 7966 : data = 8'h00;
 7967 : data = 8'h00;
 7968 : data = 8'h00;
 7969 : data = 8'h00;
 7970 : data = 8'h00;
 7971 : data = 8'h00;
 7972 : data = 8'h00;
 7973 : data = 8'h00;
 7974 : data = 8'h00;
 7975 : data = 8'h00;
 7976 : data = 8'h00;
 7977 : data = 8'h00;
 7978 : data = 8'h00;
 7979 : data = 8'h00;
 7980 : data = 8'h00;
 7981 : data = 8'h00;
 7982 : data = 8'h00;
 7983 : data = 8'h00;
 7984 : data = 8'h00;
 7985 : data = 8'h00;
 7986 : data = 8'h00;
 7987 : data = 8'h00;
 7988 : data = 8'h00;
 7989 : data = 8'h00;
 7990 : data = 8'h00;
 7991 : data = 8'h00;
 7992 : data = 8'h00;
 7993 : data = 8'h00;
 7994 : data = 8'h00;
 7995 : data = 8'h00;
 7996 : data = 8'h00;
 7997 : data = 8'h00;
 7998 : data = 8'h00;
 7999 : data = 8'h00;
 8000 : data = 8'h00;
 8001 : data = 8'h00;
 8002 : data = 8'h00;
 8003 : data = 8'h00;
 8004 : data = 8'h00;
 8005 : data = 8'h00;
 8006 : data = 8'h00;
 8007 : data = 8'h00;
 8008 : data = 8'h00;
 8009 : data = 8'h00;
 8010 : data = 8'h00;
 8011 : data = 8'h00;
 8012 : data = 8'h00;
 8013 : data = 8'h00;
 8014 : data = 8'h00;
 8015 : data = 8'h00;
 8016 : data = 8'h00;
 8017 : data = 8'h00;
 8018 : data = 8'h00;
 8019 : data = 8'h00;
 8020 : data = 8'h00;
 8021 : data = 8'h00;
 8022 : data = 8'h00;
 8023 : data = 8'h00;
 8024 : data = 8'h00;
 8025 : data = 8'h00;
 8026 : data = 8'h00;
 8027 : data = 8'h00;
 8028 : data = 8'h00;
 8029 : data = 8'h00;
 8030 : data = 8'h00;
 8031 : data = 8'h00;
 8032 : data = 8'h00;
 8033 : data = 8'h00;
 8034 : data = 8'h00;
 8035 : data = 8'h00;
 8036 : data = 8'h00;
 8037 : data = 8'h00;
 8038 : data = 8'h00;
 8039 : data = 8'h00;
 8040 : data = 8'h00;
 8041 : data = 8'h00;
 8042 : data = 8'h00;
 8043 : data = 8'h00;
 8044 : data = 8'h00;
 8045 : data = 8'h00;
 8046 : data = 8'h00;
 8047 : data = 8'h00;
 8048 : data = 8'h00;
 8049 : data = 8'h00;
 8050 : data = 8'h00;
 8051 : data = 8'h00;
 8052 : data = 8'h00;
 8053 : data = 8'h00;
 8054 : data = 8'h00;
 8055 : data = 8'h00;
 8056 : data = 8'h00;
 8057 : data = 8'h00;
 8058 : data = 8'h00;
 8059 : data = 8'h00;
 8060 : data = 8'h00;
 8061 : data = 8'h00;
 8062 : data = 8'h00;
 8063 : data = 8'h00;
 8064 : data = 8'h00;
 8065 : data = 8'h00;
 8066 : data = 8'h00;
 8067 : data = 8'h00;
 8068 : data = 8'h00;
 8069 : data = 8'h00;
 8070 : data = 8'h00;
 8071 : data = 8'h00;
 8072 : data = 8'h00;
 8073 : data = 8'h00;
 8074 : data = 8'h00;
 8075 : data = 8'h00;
 8076 : data = 8'h00;
 8077 : data = 8'h00;
 8078 : data = 8'h00;
 8079 : data = 8'h00;
 8080 : data = 8'h00;
 8081 : data = 8'h00;
 8082 : data = 8'h00;
 8083 : data = 8'h00;
 8084 : data = 8'h00;
 8085 : data = 8'h00;
 8086 : data = 8'h00;
 8087 : data = 8'h00;
 8088 : data = 8'h00;
 8089 : data = 8'h00;
 8090 : data = 8'h00;
 8091 : data = 8'h00;
 8092 : data = 8'h00;
 8093 : data = 8'h00;
 8094 : data = 8'h00;
 8095 : data = 8'h00;
 8096 : data = 8'h00;
 8097 : data = 8'h00;
 8098 : data = 8'h00;
 8099 : data = 8'h00;
 8100 : data = 8'h00;
 8101 : data = 8'h00;
 8102 : data = 8'h00;
 8103 : data = 8'h00;
 8104 : data = 8'h00;
 8105 : data = 8'h00;
 8106 : data = 8'h00;
 8107 : data = 8'h00;
 8108 : data = 8'h00;
 8109 : data = 8'h00;
 8110 : data = 8'h00;
 8111 : data = 8'h00;
 8112 : data = 8'h00;
 8113 : data = 8'h00;
 8114 : data = 8'h00;
 8115 : data = 8'h00;
 8116 : data = 8'h00;
 8117 : data = 8'h00;
 8118 : data = 8'h00;
 8119 : data = 8'h00;
 8120 : data = 8'h00;
 8121 : data = 8'h00;
 8122 : data = 8'h00;
 8123 : data = 8'h00;
 8124 : data = 8'h00;
 8125 : data = 8'h00;
 8126 : data = 8'h00;
 8127 : data = 8'h00;
 8128 : data = 8'h00;
 8129 : data = 8'h00;
 8130 : data = 8'h00;
 8131 : data = 8'h00;
 8132 : data = 8'h00;
 8133 : data = 8'h00;
 8134 : data = 8'h00;
 8135 : data = 8'h00;
 8136 : data = 8'h00;
 8137 : data = 8'h00;
 8138 : data = 8'h00;
 8139 : data = 8'h00;
 8140 : data = 8'h00;
 8141 : data = 8'h00;
 8142 : data = 8'h00;
 8143 : data = 8'h00;
 8144 : data = 8'h00;
 8145 : data = 8'h00;
 8146 : data = 8'h00;
 8147 : data = 8'h00;
 8148 : data = 8'h00;
 8149 : data = 8'h00;
 8150 : data = 8'h00;
 8151 : data = 8'h00;
 8152 : data = 8'h00;
 8153 : data = 8'h00;
 8154 : data = 8'h00;
 8155 : data = 8'h00;
 8156 : data = 8'h00;
 8157 : data = 8'h00;
 8158 : data = 8'h00;
 8159 : data = 8'h00;
 8160 : data = 8'h00;
 8161 : data = 8'h00;
 8162 : data = 8'h00;
 8163 : data = 8'h00;
 8164 : data = 8'h00;
 8165 : data = 8'h00;
 8166 : data = 8'h00;
 8167 : data = 8'h00;
 8168 : data = 8'h00;
 8169 : data = 8'h00;
 8170 : data = 8'h00;
 8171 : data = 8'h00;
 8172 : data = 8'h00;
 8173 : data = 8'h00;
 8174 : data = 8'h00;
 8175 : data = 8'h00;
 8176 : data = 8'h00;
 8177 : data = 8'h00;
 8178 : data = 8'h00;
 8179 : data = 8'h00;
 8180 : data = 8'h00;
 8181 : data = 8'h00;
 8182 : data = 8'h00;
 8183 : data = 8'h00;
 8184 : data = 8'h00;
 8185 : data = 8'h00;
 8186 : data = 8'h00;
 8187 : data = 8'h00;
 8188 : data = 8'h00;
 8189 : data = 8'h00;
 8190 : data = 8'h00;
 8191 : data = 8'h00;
 8192 : data = 8'hFF;
 8193 : data = 8'hFF;
 8194 : data = 8'hFF;
 8195 : data = 8'hFF;
 8196 : data = 8'hFF;
 8197 : data = 8'hFF;
 8198 : data = 8'hFF;
 8199 : data = 8'hFF;
 8200 : data = 8'hFF;
 8201 : data = 8'hFF;
 8202 : data = 8'hFF;
 8203 : data = 8'hFF;
 8204 : data = 8'hFF;
 8205 : data = 8'hFF;
 8206 : data = 8'hFF;
 8207 : data = 8'hFF;
 8208 : data = 8'hFF;
 8209 : data = 8'hFF;
 8210 : data = 8'hFF;
 8211 : data = 8'hFF;
 8212 : data = 8'hFF;
 8213 : data = 8'hFF;
 8214 : data = 8'hFF;
 8215 : data = 8'hFF;
 8216 : data = 8'hFF;
 8217 : data = 8'hFF;
 8218 : data = 8'hFF;
 8219 : data = 8'hFF;
 8220 : data = 8'hFF;
 8221 : data = 8'hFF;
 8222 : data = 8'hFF;
 8223 : data = 8'hFF;
 8224 : data = 8'hFF;
 8225 : data = 8'hFF;
 8226 : data = 8'hFF;
 8227 : data = 8'hFF;
 8228 : data = 8'hFF;
 8229 : data = 8'hFF;
 8230 : data = 8'hFF;
 8231 : data = 8'hFF;
 8232 : data = 8'hFF;
 8233 : data = 8'hFF;
 8234 : data = 8'hFF;
 8235 : data = 8'hFF;
 8236 : data = 8'hFF;
 8237 : data = 8'hFF;
 8238 : data = 8'hFF;
 8239 : data = 8'hFF;
 8240 : data = 8'hFF;
 8241 : data = 8'hFF;
 8242 : data = 8'hFF;
 8243 : data = 8'hFF;
 8244 : data = 8'hFF;
 8245 : data = 8'hFF;
 8246 : data = 8'hFF;
 8247 : data = 8'hFF;
 8248 : data = 8'hFF;
 8249 : data = 8'hFF;
 8250 : data = 8'hFF;
 8251 : data = 8'hFF;
 8252 : data = 8'hFF;
 8253 : data = 8'hFF;
 8254 : data = 8'hFF;
 8255 : data = 8'hFF;
 8256 : data = 8'hFF;
 8257 : data = 8'hFF;
 8258 : data = 8'hFF;
 8259 : data = 8'hFF;
 8260 : data = 8'hFF;
 8261 : data = 8'hFF;
 8262 : data = 8'hFF;
 8263 : data = 8'hFF;
 8264 : data = 8'hFF;
 8265 : data = 8'hFF;
 8266 : data = 8'hFF;
 8267 : data = 8'hFF;
 8268 : data = 8'hFF;
 8269 : data = 8'hFF;
 8270 : data = 8'hFF;
 8271 : data = 8'hFF;
 8272 : data = 8'hFF;
 8273 : data = 8'hFF;
 8274 : data = 8'hFF;
 8275 : data = 8'hFF;
 8276 : data = 8'hFF;
 8277 : data = 8'hFF;
 8278 : data = 8'hFF;
 8279 : data = 8'hFF;
 8280 : data = 8'hFF;
 8281 : data = 8'hFF;
 8282 : data = 8'hFF;
 8283 : data = 8'hFF;
 8284 : data = 8'hFF;
 8285 : data = 8'hFF;
 8286 : data = 8'hFF;
 8287 : data = 8'hFF;
 8288 : data = 8'hFF;
 8289 : data = 8'hFF;
 8290 : data = 8'hFF;
 8291 : data = 8'hFF;
 8292 : data = 8'h00;
 8293 : data = 8'h00;
 8294 : data = 8'h00;
 8295 : data = 8'h00;
 8296 : data = 8'h00;
 8297 : data = 8'h00;
 8298 : data = 8'h00;
 8299 : data = 8'h00;
 8300 : data = 8'h00;
 8301 : data = 8'h00;
 8302 : data = 8'h00;
 8303 : data = 8'h00;
 8304 : data = 8'h00;
 8305 : data = 8'h00;
 8306 : data = 8'h00;
 8307 : data = 8'h00;
 8308 : data = 8'h00;
 8309 : data = 8'h00;
 8310 : data = 8'h00;
 8311 : data = 8'h00;
 8312 : data = 8'h00;
 8313 : data = 8'h00;
 8314 : data = 8'h00;
 8315 : data = 8'h00;
 8316 : data = 8'h00;
 8317 : data = 8'h00;
 8318 : data = 8'h00;
 8319 : data = 8'h00;
 8320 : data = 8'h00;
 8321 : data = 8'h00;
 8322 : data = 8'h00;
 8323 : data = 8'h00;
 8324 : data = 8'h00;
 8325 : data = 8'h00;
 8326 : data = 8'h00;
 8327 : data = 8'h00;
 8328 : data = 8'h00;
 8329 : data = 8'h00;
 8330 : data = 8'h00;
 8331 : data = 8'h00;
 8332 : data = 8'h00;
 8333 : data = 8'h00;
 8334 : data = 8'h00;
 8335 : data = 8'h00;
 8336 : data = 8'h00;
 8337 : data = 8'h00;
 8338 : data = 8'h00;
 8339 : data = 8'h00;
 8340 : data = 8'h00;
 8341 : data = 8'h00;
 8342 : data = 8'h00;
 8343 : data = 8'h00;
 8344 : data = 8'h00;
 8345 : data = 8'h00;
 8346 : data = 8'h00;
 8347 : data = 8'h00;
 8348 : data = 8'h00;
 8349 : data = 8'h00;
 8350 : data = 8'h00;
 8351 : data = 8'h00;
 8352 : data = 8'h00;
 8353 : data = 8'h00;
 8354 : data = 8'h00;
 8355 : data = 8'h00;
 8356 : data = 8'h00;
 8357 : data = 8'h00;
 8358 : data = 8'h00;
 8359 : data = 8'h00;
 8360 : data = 8'h00;
 8361 : data = 8'h00;
 8362 : data = 8'h00;
 8363 : data = 8'h00;
 8364 : data = 8'h00;
 8365 : data = 8'h00;
 8366 : data = 8'h00;
 8367 : data = 8'h00;
 8368 : data = 8'h00;
 8369 : data = 8'h00;
 8370 : data = 8'h00;
 8371 : data = 8'h00;
 8372 : data = 8'h00;
 8373 : data = 8'h00;
 8374 : data = 8'h00;
 8375 : data = 8'h00;
 8376 : data = 8'h00;
 8377 : data = 8'h00;
 8378 : data = 8'h00;
 8379 : data = 8'h00;
 8380 : data = 8'h00;
 8381 : data = 8'h00;
 8382 : data = 8'h00;
 8383 : data = 8'h00;
 8384 : data = 8'h00;
 8385 : data = 8'h00;
 8386 : data = 8'h00;
 8387 : data = 8'h00;
 8388 : data = 8'h00;
 8389 : data = 8'h00;
 8390 : data = 8'h00;
 8391 : data = 8'h00;
 8392 : data = 8'h00;
 8393 : data = 8'h00;
 8394 : data = 8'h00;
 8395 : data = 8'h00;
 8396 : data = 8'h00;
 8397 : data = 8'h00;
 8398 : data = 8'h00;
 8399 : data = 8'h00;
 8400 : data = 8'h00;
 8401 : data = 8'h00;
 8402 : data = 8'h00;
 8403 : data = 8'h00;
 8404 : data = 8'h00;
 8405 : data = 8'h00;
 8406 : data = 8'h00;
 8407 : data = 8'h00;
 8408 : data = 8'h00;
 8409 : data = 8'h00;
 8410 : data = 8'h00;
 8411 : data = 8'h00;
 8412 : data = 8'h00;
 8413 : data = 8'h00;
 8414 : data = 8'h00;
 8415 : data = 8'h00;
 8416 : data = 8'h00;
 8417 : data = 8'h00;
 8418 : data = 8'h00;
 8419 : data = 8'h00;
 8420 : data = 8'h00;
 8421 : data = 8'h00;
 8422 : data = 8'h00;
 8423 : data = 8'h00;
 8424 : data = 8'h00;
 8425 : data = 8'h00;
 8426 : data = 8'h00;
 8427 : data = 8'h00;
 8428 : data = 8'h00;
 8429 : data = 8'h00;
 8430 : data = 8'h00;
 8431 : data = 8'h00;
 8432 : data = 8'h00;
 8433 : data = 8'h00;
 8434 : data = 8'h00;
 8435 : data = 8'h00;
 8436 : data = 8'h00;
 8437 : data = 8'h00;
 8438 : data = 8'h00;
 8439 : data = 8'h00;
 8440 : data = 8'h00;
 8441 : data = 8'h00;
 8442 : data = 8'h00;
 8443 : data = 8'h00;
 8444 : data = 8'h00;
 8445 : data = 8'h00;
 8446 : data = 8'h00;
 8447 : data = 8'h00;
 8448 : data = 8'h80;
 8449 : data = 8'h00;
 8450 : data = 8'h00;
 8451 : data = 8'h00;
 8452 : data = 8'h00;
 8453 : data = 8'h00;
 8454 : data = 8'h00;
 8455 : data = 8'h00;
 8456 : data = 8'h00;
 8457 : data = 8'h00;
 8458 : data = 8'h00;
 8459 : data = 8'h00;
 8460 : data = 8'h00;
 8461 : data = 8'h00;
 8462 : data = 8'h00;
 8463 : data = 8'h00;
 8464 : data = 8'h00;
 8465 : data = 8'h00;
 8466 : data = 8'h00;
 8467 : data = 8'h00;
 8468 : data = 8'h00;
 8469 : data = 8'h00;
 8470 : data = 8'h00;
 8471 : data = 8'h00;
 8472 : data = 8'h00;
 8473 : data = 8'h00;
 8474 : data = 8'h00;
 8475 : data = 8'h00;
 8476 : data = 8'h00;
 8477 : data = 8'h00;
 8478 : data = 8'h00;
 8479 : data = 8'h00;
 8480 : data = 8'h00;
 8481 : data = 8'h00;
 8482 : data = 8'h00;
 8483 : data = 8'h00;
 8484 : data = 8'h00;
 8485 : data = 8'h00;
 8486 : data = 8'h00;
 8487 : data = 8'h00;
 8488 : data = 8'h00;
 8489 : data = 8'h00;
 8490 : data = 8'h00;
 8491 : data = 8'h00;
 8492 : data = 8'h00;
 8493 : data = 8'h00;
 8494 : data = 8'h00;
 8495 : data = 8'h00;
 8496 : data = 8'h00;
 8497 : data = 8'h00;
 8498 : data = 8'h00;
 8499 : data = 8'h00;
 8500 : data = 8'h00;
 8501 : data = 8'h00;
 8502 : data = 8'h00;
 8503 : data = 8'h00;
 8504 : data = 8'h00;
 8505 : data = 8'h00;
 8506 : data = 8'h00;
 8507 : data = 8'h00;
 8508 : data = 8'h00;
 8509 : data = 8'h00;
 8510 : data = 8'h00;
 8511 : data = 8'h00;
 8512 : data = 8'h00;
 8513 : data = 8'h00;
 8514 : data = 8'h00;
 8515 : data = 8'h00;
 8516 : data = 8'h00;
 8517 : data = 8'h00;
 8518 : data = 8'h00;
 8519 : data = 8'h00;
 8520 : data = 8'h00;
 8521 : data = 8'h00;
 8522 : data = 8'h00;
 8523 : data = 8'h00;
 8524 : data = 8'h00;
 8525 : data = 8'h00;
 8526 : data = 8'h00;
 8527 : data = 8'h00;
 8528 : data = 8'h00;
 8529 : data = 8'h00;
 8530 : data = 8'h00;
 8531 : data = 8'h00;
 8532 : data = 8'h00;
 8533 : data = 8'h00;
 8534 : data = 8'h00;
 8535 : data = 8'h00;
 8536 : data = 8'h00;
 8537 : data = 8'h00;
 8538 : data = 8'h00;
 8539 : data = 8'h00;
 8540 : data = 8'h00;
 8541 : data = 8'h00;
 8542 : data = 8'h00;
 8543 : data = 8'h00;
 8544 : data = 8'h00;
 8545 : data = 8'h00;
 8546 : data = 8'h00;
 8547 : data = 8'h00;
 8548 : data = 8'h00;
 8549 : data = 8'h00;
 8550 : data = 8'h00;
 8551 : data = 8'h00;
 8552 : data = 8'h00;
 8553 : data = 8'h00;
 8554 : data = 8'h00;
 8555 : data = 8'h00;
 8556 : data = 8'h00;
 8557 : data = 8'h00;
 8558 : data = 8'h00;
 8559 : data = 8'h00;
 8560 : data = 8'h00;
 8561 : data = 8'h00;
 8562 : data = 8'h00;
 8563 : data = 8'h00;
 8564 : data = 8'h00;
 8565 : data = 8'h00;
 8566 : data = 8'h00;
 8567 : data = 8'h00;
 8568 : data = 8'h00;
 8569 : data = 8'h00;
 8570 : data = 8'h00;
 8571 : data = 8'h00;
 8572 : data = 8'h00;
 8573 : data = 8'h00;
 8574 : data = 8'h00;
 8575 : data = 8'h00;
 8576 : data = 8'h00;
 8577 : data = 8'h00;
 8578 : data = 8'h00;
 8579 : data = 8'h00;
 8580 : data = 8'h00;
 8581 : data = 8'h00;
 8582 : data = 8'h00;
 8583 : data = 8'h00;
 8584 : data = 8'h00;
 8585 : data = 8'h00;
 8586 : data = 8'h00;
 8587 : data = 8'h00;
 8588 : data = 8'h00;
 8589 : data = 8'h00;
 8590 : data = 8'h00;
 8591 : data = 8'h00;
 8592 : data = 8'h00;
 8593 : data = 8'h00;
 8594 : data = 8'h00;
 8595 : data = 8'h00;
 8596 : data = 8'h00;
 8597 : data = 8'h00;
 8598 : data = 8'h00;
 8599 : data = 8'h00;
 8600 : data = 8'h00;
 8601 : data = 8'h00;
 8602 : data = 8'h00;
 8603 : data = 8'h00;
 8604 : data = 8'h00;
 8605 : data = 8'h00;
 8606 : data = 8'h00;
 8607 : data = 8'h00;
 8608 : data = 8'h00;
 8609 : data = 8'h00;
 8610 : data = 8'h00;
 8611 : data = 8'h00;
 8612 : data = 8'h00;
 8613 : data = 8'h00;
 8614 : data = 8'h00;
 8615 : data = 8'h00;
 8616 : data = 8'h00;
 8617 : data = 8'h00;
 8618 : data = 8'h00;
 8619 : data = 8'h00;
 8620 : data = 8'h00;
 8621 : data = 8'h00;
 8622 : data = 8'h00;
 8623 : data = 8'h00;
 8624 : data = 8'h00;
 8625 : data = 8'h00;
 8626 : data = 8'h00;
 8627 : data = 8'h00;
 8628 : data = 8'h00;
 8629 : data = 8'h00;
 8630 : data = 8'h00;
 8631 : data = 8'h00;
 8632 : data = 8'h00;
 8633 : data = 8'h00;
 8634 : data = 8'h00;
 8635 : data = 8'h00;
 8636 : data = 8'h00;
 8637 : data = 8'h00;
 8638 : data = 8'h00;
 8639 : data = 8'h00;
 8640 : data = 8'h00;
 8641 : data = 8'h00;
 8642 : data = 8'h00;
 8643 : data = 8'h00;
 8644 : data = 8'h00;
 8645 : data = 8'h00;
 8646 : data = 8'h00;
 8647 : data = 8'h00;
 8648 : data = 8'h00;
 8649 : data = 8'h00;
 8650 : data = 8'h00;
 8651 : data = 8'h00;
 8652 : data = 8'h00;
 8653 : data = 8'h00;
 8654 : data = 8'h00;
 8655 : data = 8'h00;
 8656 : data = 8'h00;
 8657 : data = 8'h00;
 8658 : data = 8'h00;
 8659 : data = 8'h00;
 8660 : data = 8'h00;
 8661 : data = 8'h00;
 8662 : data = 8'h00;
 8663 : data = 8'h00;
 8664 : data = 8'h00;
 8665 : data = 8'h00;
 8666 : data = 8'h00;
 8667 : data = 8'h00;
 8668 : data = 8'h00;
 8669 : data = 8'h00;
 8670 : data = 8'h00;
 8671 : data = 8'h00;
 8672 : data = 8'h00;
 8673 : data = 8'h00;
 8674 : data = 8'h00;
 8675 : data = 8'h00;
 8676 : data = 8'h00;
 8677 : data = 8'h00;
 8678 : data = 8'h00;
 8679 : data = 8'h00;
 8680 : data = 8'h00;
 8681 : data = 8'h00;
 8682 : data = 8'h00;
 8683 : data = 8'h00;
 8684 : data = 8'h00;
 8685 : data = 8'h00;
 8686 : data = 8'h00;
 8687 : data = 8'h00;
 8688 : data = 8'h00;
 8689 : data = 8'h00;
 8690 : data = 8'h00;
 8691 : data = 8'h00;
 8692 : data = 8'h00;
 8693 : data = 8'h00;
 8694 : data = 8'h00;
 8695 : data = 8'h00;
 8696 : data = 8'h00;
 8697 : data = 8'h00;
 8698 : data = 8'h00;
 8699 : data = 8'h00;
 8700 : data = 8'h00;
 8701 : data = 8'h00;
 8702 : data = 8'h00;
 8703 : data = 8'h00;
 8704 : data = 8'h04;
 8705 : data = 8'h00;
 8706 : data = 8'h00;
 8707 : data = 8'h00;
 default: data = 8'h01; // invalid instruction
 endcase
end
endmodule
